-- GENERATED WITH MATLAB...

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package CE_5G_pkg is 


type type_m291a2int is array (0 to 290,0 to 1) of integer range 0 to 3; 
type type_m4a2x16std is array (0 to 4-1,0 to 2-1) of std_logic_vector(16-1 downto 0); 

constant dict_DMRS : type_m4a2x16std := ( 
 	 ("1010010101111101","1010010101111101"), 
  	 ("0101101010000011","1010010101111101"), 
  	 ("0101101010000011","0101101010000011"), 
  	 ("1010010101111101","0101101010000011")); 

constant dictInd_DMRS : type_m291a2int := ( 
	 (1,1), 
	 (3,0), 
	 (1,1), 
	 (2,1), 
	 (2,3), 
	 (0,1), 
	 (1,1), 
	 (1,1), 
	 (0,0), 
	 (3,1), 
	 (3,1), 
	 (2,2), 
	 (0,1), 
	 (0,0), 
	 (1,3), 
	 (2,2), 
	 (3,3), 
	 (0,0), 
	 (1,2), 
	 (2,2), 
	 (3,2), 
	 (0,2), 
	 (0,0), 
	 (2,1), 
	 (0,3), 
	 (2,3), 
	 (0,3), 
	 (2,0), 
	 (3,2), 
	 (1,3), 
	 (3,0), 
	 (0,2), 
	 (2,0), 
	 (1,1), 
	 (0,1), 
	 (0,0), 
	 (3,3), 
	 (3,0), 
	 (3,2), 
	 (1,3), 
	 (1,2), 
	 (3,0), 
	 (2,3), 
	 (1,0), 
	 (1,1), 
	 (2,1), 
	 (1,0), 
	 (2,1), 
	 (3,0), 
	 (0,2), 
	 (0,3), 
	 (2,2), 
	 (3,2), 
	 (3,3), 
	 (1,1), 
	 (2,3), 
	 (2,2), 
	 (1,2), 
	 (0,1), 
	 (2,0), 
	 (3,1), 
	 (0,1), 
	 (2,3), 
	 (0,0), 
	 (0,3), 
	 (0,1), 
	 (2,1), 
	 (3,0), 
	 (2,2), 
	 (1,3), 
	 (2,1), 
	 (1,1), 
	 (3,2), 
	 (2,2), 
	 (1,2), 
	 (2,1), 
	 (2,0), 
	 (0,3), 
	 (3,2), 
	 (0,3), 
	 (1,0), 
	 (1,2), 
	 (0,3), 
	 (1,0), 
	 (1,0), 
	 (1,0), 
	 (1,3), 
	 (2,3), 
	 (3,3), 
	 (3,2), 
	 (0,0), 
	 (0,2), 
	 (1,2), 
	 (2,2), 
	 (1,2), 
	 (3,0), 
	 (0,1), 
	 (3,1), 
	 (1,0), 
	 (3,1), 
	 (3,0), 
	 (2,3), 
	 (2,0), 
	 (3,2), 
	 (0,1), 
	 (2,3), 
	 (2,3), 
	 (1,3), 
	 (3,2), 
	 (3,2), 
	 (3,2), 
	 (2,2), 
	 (0,1), 
	 (2,1), 
	 (3,0), 
	 (2,0), 
	 (2,1), 
	 (0,2), 
	 (3,2), 
	 (3,2), 
	 (2,3), 
	 (1,3), 
	 (1,1), 
	 (1,3), 
	 (2,0), 
	 (2,3), 
	 (1,2), 
	 (0,3), 
	 (0,1), 
	 (1,0), 
	 (1,0), 
	 (2,0), 
	 (1,2), 
	 (2,1), 
	 (2,0), 
	 (3,2), 
	 (1,3), 
	 (3,3), 
	 (0,1), 
	 (2,2), 
	 (2,3), 
	 (2,3), 
	 (2,3), 
	 (2,1), 
	 (0,1), 
	 (2,2), 
	 (2,0), 
	 (3,1), 
	 (0,2), 
	 (1,0), 
	 (0,2), 
	 (2,3), 
	 (2,0), 
	 (1,0), 
	 (1,0), 
	 (3,0), 
	 (3,2), 
	 (3,1), 
	 (1,3), 
	 (3,0), 
	 (2,3), 
	 (1,1), 
	 (1,0), 
	 (3,2), 
	 (1,2), 
	 (3,3), 
	 (0,2), 
	 (1,2), 
	 (2,1), 
	 (0,1), 
	 (3,3), 
	 (0,2), 
	 (3,3), 
	 (3,0), 
	 (3,3), 
	 (2,0), 
	 (1,2), 
	 (2,3), 
	 (3,3), 
	 (1,0), 
	 (3,1), 
	 (0,0), 
	 (1,1), 
	 (3,2), 
	 (0,3), 
	 (1,1), 
	 (0,2), 
	 (2,1), 
	 (0,0), 
	 (0,3), 
	 (3,1), 
	 (0,3), 
	 (1,0), 
	 (3,0), 
	 (0,2), 
	 (0,3), 
	 (0,0), 
	 (1,2), 
	 (3,3), 
	 (1,2), 
	 (2,3), 
	 (0,0), 
	 (3,2), 
	 (0,0), 
	 (1,2), 
	 (0,2), 
	 (3,3), 
	 (0,3), 
	 (2,0), 
	 (0,0), 
	 (1,0), 
	 (0,1), 
	 (2,1), 
	 (0,0), 
	 (3,3), 
	 (2,0), 
	 (2,0), 
	 (0,1), 
	 (2,0), 
	 (0,2), 
	 (1,3), 
	 (1,3), 
	 (3,0), 
	 (3,3), 
	 (1,1), 
	 (3,3), 
	 (3,3), 
	 (2,3), 
	 (0,3), 
	 (1,3), 
	 (1,1), 
	 (3,0), 
	 (2,0), 
	 (1,3), 
	 (3,3), 
	 (0,3), 
	 (3,2), 
	 (0,2), 
	 (1,3), 
	 (2,2), 
	 (3,2), 
	 (3,0), 
	 (0,0), 
	 (3,3), 
	 (0,1), 
	 (1,3), 
	 (1,2), 
	 (3,3), 
	 (3,2), 
	 (0,1), 
	 (0,1), 
	 (3,2), 
	 (3,1), 
	 (0,1), 
	 (3,0), 
	 (1,3), 
	 (0,2), 
	 (1,1), 
	 (3,1), 
	 (1,2), 
	 (1,2), 
	 (2,0), 
	 (1,0), 
	 (3,1), 
	 (1,1), 
	 (1,3), 
	 (3,2), 
	 (2,3), 
	 (0,0), 
	 (0,2), 
	 (3,1), 
	 (2,3), 
	 (2,1), 
	 (0,2), 
	 (1,0), 
	 (2,0), 
	 (3,2), 
	 (1,3), 
	 (1,3), 
	 (2,2), 
	 (0,1), 
	 (0,1), 
	 (0,0), 
	 (1,3), 
	 (3,3), 
	 (2,2), 
	 (1,2), 
	 (2,0), 
	 (2,0), 
	 (2,1), 
	 (2,1)); 

end CE_5G_pkg; 
