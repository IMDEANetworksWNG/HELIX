

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
giSbz6lFREHMEDzBP8fkL+cjyMAzxx4373IBs3k0mBF0lyQV5MR794C4py6ITwcsR6aK++Utvfz3
Z9Wb2XVKWg==


`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
OHsjOqigLPnUdhYo4s7q/8keAnfBnTUsSx0jR3kWaBW7MFMEBGz4ilTIx67/xkyzJSWMNFxgcNeo
NYflRvGJBfMgj+mOhl4K/rSvdLy0PYQqaIBKtW3r3bYyIoM0vfYjAhgRNG5+CyFjqoCTGLp5J0BO
AAn93ce3Ri/CgHnSt3c=


`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
YGiXz7o4JhofQ0AokPo7aVVC5313FmyTmDeXZpQmTdhCCABBeFTpwucOcjjw3bDkubDhzLfDro3/
s+btR6bljbMKeOykv04xCACdlAScehaiNLcGgTM7IWDwiReb+FJs3plZAC8VTisbXHOqQad/6CWW
KXAb/G/DLL1LPbpabHO/Ky6yeXFp4CX1Z0sprGf97cbBc7nqJkYr2xzism1SDnGGw7yTez5Jg3xP
NsZXePlctk8FOEkov6/seR8xVFtOM8p360/ktKBqgpDrBesIiggmYqlD3NQ7EqAhSDOVhHziPub0
DQEyku9jztTFEKSAEwiwi9Qv3k5HHBkjIzkCyg==


`pragma protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KGrUMg5ySDiN3C2YRpbBsg7x76hfgEpVeEWSihjwXT3R+wiFbM68xaw5yHG7YwMeiYg3+Rw9Z/Oy
mcsGg8uaRLn2rUElUYaFvkpHEkqgh36ESByM2Ux75jAL5HMT7vue1YNiekQbtkK+7cmbcGbYFF11
945Y0rY8L5YeDgUUheXw9AqZaz/0K5/GHGQCeiDhP9EW2cCaesuuwi3xDQzNRsKUshLwwhzxnjwe
TsHjw0FF69ZkYNgVJY4xHy1Z2/STXr/bRp8i0x4nW9EvPoUR+NmV5Y1KpHeSqy+GaWDre32c2re6
0Ps6wCWy8nKhhLsSYQQLe+vpTHKyYH9mWU3+ww==


`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
cPHrJ+aktiD6VmpJxfzG17f5ApguZrVZ+hoAdVfqMzBI4Bf7miweJPMHQAP3lm5F4DJpvHkD5U1c
1yCklGy4KC1aEslOOJdRrNW7iraFNmRIoKkbUX0j4cWUT8XhQil9uGGNb7ah3ZGla1HC5SoviUHZ
CPHWnj1Ex+dEStvjyfV5sozPqRmGgv6pDe1BDzj3Gn9sgCEKhAW82x4Ms6J702gKUnzkuvtqQcq6
gJHcYmvG/7f681rZr7sSdcZU2XU7cNWOFnJoXlP5gODD4yPvAgs2RXco/s8qwED8LpesYJce6Y5t
Gy1JOhE6wynPObsiIK1ivg+5AaHqReh0x+ojjQ==


`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
knEP1CoC7G1uOBV6pcAuqxmxi8zefOeS7D+f8C1AlyJ5Peux0yDrKfej7ZfbHNTlslsz57imA6mT
6OlpXnmMKl2/saV8eOjMopAct4XrV+9Rpw9PEunNOeMgZpaPA+bf81ZRAkdBSC/UwHBZ18z+2Sef
NXANmK6nWz5OxDpQ4LQ=


`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OewN470bZRWGUqHttYxO5MD4x67TksEKsV4DP0z015Xd4FzLVfsuapLLsHZvm7xXCLSbnPt62ijo
1kxLS/9MQDo2lhw+aj86bjyBAZbmC/ihnH4phAkM3ah9lLrx4GsaMeGZcllOxhtnB/0BccDmTXMM
gaHcfeaM7bsFB7BI0koMCOx7YtMreR3jaHLo5ZDI43/0rXFQuEMxqCBBM6dieaJ9AAonkrNNjMhY
s0+OsAoTJXdyHGw/Z7RndEfKqoF0ocyprizehXKKCHeXAyvw1NxiOwEuRd/bWUu0KOtcJdIkhZQY
Q2BQrm8YhOfEdVGMowquIwxA3m8rybWjkOUQEA==


`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 479680)
`pragma protect data_block
se3q5e3u3ZpNDq3isdundILs7UQRSZsweTcLaa3IBkUuwh8r79Rj2n1kZ6KjL9Ks7Zk+szu2UTzI
NPBnGeJvwuJDBfux5+xWYKQ/sJfyefOVRYXtr7IckhFZsoztnw6RBLJV7hX4QG4lYoBsDmSLJQFg
u3cPZXqtN3h3XZj5SlCsJEs328/fW4GSVw5x9GV6p16mvVZYiAfEURris/72A0Njo6pBrLDoB60/
nN8Ax3cYnI2WCXpFWfkmZiYavGaIwQKt4L+zOXq4ocbcwOTxrjZLWI1kC1mbplEJXc0Qw2jfHqy3
3yYsJ3amJwQT0jA/C0pjJ+pN1ab9KS0yNCWyMRif4ykjyXbFpvHNx18U9XdidJPSRT70sgTFV89N
6LTMwBFPhL2TJ9eVKOTKlN24UAIB9QbCAjRsTXkA1myB/4X08kldodOyV9wAWrhro3GG2Cq7u4bh
VTm8D58/VNcFJ6TvpKT/it5U0T71FigxI5piiFiRUQO0abNOi4qLSSyak5e/5DYyQ1XkwW+FPx3N
dbvOFAvUidAp2WbIpYbBuyZV0O9Gcdv1+3zOAWE9vMokqauPxHPbxfzRRfTjfJflcl8yfB08xVMy
v/7wjJCrr3wxEJwR2SN2u8vSQkMzvkvkU0lGYj5Kpn0v6CZ3iBBFCzm1MgRON+whmEww3anpRanN
PUiEjPCH2ORJ1Y4faKugUdkLQosXy0VJ6h7t5Gxpk/Te1mbXOWMl3XMEX6ErXY5sOVD1/l0FimU6
/rBq56IIXGwdec/4QXE0ahwYc1DE27DzqDf4N3NhoPqkc9mIL/GXdzuRFtR8ogDitU3JMv3dXw2z
H/8KCbA1kcw/OuEq7iy4Wyc5mSTjOe+yFnclMYUjZVA0JzQvxa0GIfX/ET5Xn1L+Jsbw443NlOYp
RbQy4LUnr5c+onu6ym8/NmiZH9ZNvGup0Mj30JABScomABWnB9zRf8lvcVRZmgSltK85rCMWorFd
JvQgU2wlacHDYCQ56dRRrqbaIqLy1MFKDBmBYnJ8gJWRYKltUWUdUyRTbA+SHWTFUlfI0zTpImUu
0WelhsvC++15RH835R7rtKd2CN2ttMprwmonDdPQDy9StsrI8UM9SzvV2+BQO3icGXUJHWMHmdhY
fdTckL+v2sWFK1QCa68Jf50ON3KkwGdRd/KmaqTFc2kGYTIJW2cf9S0GdQQcVP31BZKI9b8KXDHR
Dz6poRbMVIC90NO/8LyLkh+DBwP48KtiZo4k306BvDtl3Bp2F6vu+f90B7VDuAc20UPDUYC8DcKt
L1Ec4oJE6+OdB5ykpma7qUqsV9OI8FeHlQxPLwv4Dz0hEiHR1eu6hyGtmSQE9NXpGRNs+sljigj5
Hw2M6Hr7SJTboGt+A1KLt7djUOO6znH9XVfW7w1QExW6HjVjZ/R4Gf1vhfDLWV6ESSK+QwqHmOY/
QFgeJfz1xPqxscl4/RNZ+UsyryUO6u6Vvyr9cjp+9omd91ScXVMp/1zWv3bq6R+wpVgrKU93B17H
04RTeFTjCMUFqOaujPZe1mqnSnMTPNQTzokKNXsZNO4S1F8IpkrYS7+g/Pa7h6YGlvKalGwfjo5D
7Bn5VYyqMN8XNJ+LspjIlLmRb0/bjbWjfyJiWO58vf7XxifhXjaoGEPOvHyRawAr3U78EB73FPl8
8oQSL3L6+MKPUUVssrPBvdJl3zDT7oni4C1pSGnam0dZjcMkNisVbmTlFAC3Qmt8zacS8w1S/Qsm
1iLnzrF4JUafFCb9OUxLiX4nioSDs9zjsQ6zum+OUpvmVudWATIJpzRFj1cEjnu9V1xsq+TUOWPe
XetsXltDckfOFziSkJc3wESbsYJ7Z7beeCfqIKz2UCULmhuSUkC404hmaAnHcJvrESo7GQdASgRw
VxUTCzrqn/nbzXC2kDxHa37r5PYAiRESZFLLu/1c8BRNGNV7KBHI6HQlOrvV+FAfcMFQuo2dvShv
4CX0pgBr3XiOjg2BvzFHiOb6wbiomAVw7gYqfHi+fVitgntlEKpoQYkUGFqA/QW7QD5kQsUdzMwQ
JkRug31AlxK/iDAESdhpiWpLwmpKUPUylvC1M81n5UayRNuYKjVoUKWQ3ZyY8j5EOeLNCyOdLyrr
CGkY4812UsOquhqy5eE45IA3HFrmedt9RiFI5IyxWTlPFwa0WaNZBxKoKs8B3Hl/Lj9Nc9euct0s
Onn4alYRGNhe7nJboAu519OBkQFdegJ9OoDC9ZF7d8YZZj0Vm51sWYYbFO5tVAYHPWwleXADn+ei
e2ctDVyXdRChOMKWdncgNmLLzfp4yRZPftgVOXg/UsVvNz2gVnNqs4nmd6Gjcwy4o1lwvGjFmFF/
iTwjI9FZF8rI1fp+5MoUbC7SLlguKWD/XaSW1iBnMKTmhGB/sgCpXKIrDD3Q+kZ0ZrNv9Q8KUqwV
IcYADS97JObrHezp3odH04PTsSizitg+XS/EBs1bBdZ7Cxe15VSju1T8hm4n+sUTuARSgs8TpiuS
VfYPRdEHDcKzYP23+RCDTCTmIj9oLOB2TFYsS1xcIc+gRH59wYilsNlfgN3qCBTvPSancrt546jP
PnCCcmuE32Cb0cIz88duE4rTpW458zJiBRcZMBuG6xHySUiHkFnDyMaiCQaS7nxo4JmCzOZRqdx3
aQvqtpMpqPWMtF8qvfbsn+4mCFQQrNqpezkSJLsTU5SzFnpP4RCuxxgx46lbAt5B+sHPgQ0qZGA3
ibj8ArWjoDqs41143R7XJwU2uOE42VGjp7uzWMd0vNTWOhUz/eRHagUhOl1jhojeaX07rrcNZZwG
q9G+G2Os0ILyRvPTTFAq3b33/L/EC9X1RYgg1PWOgrwld5brbsMyYWIbGPMVRQiFEUFuDu3+JFe5
efFWYaYw4QtUeSPV9jUNJOtX8CBrq1xusf4byESznz3SPcBjoMp4xNu47nmp23PXE8IKOlCWxWvK
VJJIfriQvAiGmgO417WT73O8kIKUbgCUwIGsjumwBo/v/LYH2SpKILdYIXpfE3bCjTh/Fd9OK3RX
CMtAtGlS1z7bXXOJfsR0Hh23slNZy7evMwhErycWqItSNTXrbCpEWXImionclcQdBwURm7S9GFZI
pX+uZIHLG9EgyY7703ZLxmdqmnnmyJvjQglNKlgvsERQxaBpllpg72aE9qblkuL9SSd2meYnatpU
UTApjfLKCJQrlGJpjyEeViS5vSCkDtjBfWdUonjqBahlfvyc1CnX4A/s4Zrg9HxJ5AVZiIQkvJHW
loL0SIje5WviJpwLr+Rkl6wEwt998x3jPkEhKx6skmf63lcP7hdePQuJx5YGX3nt7xhaSxcdKpTA
C8v9p/yGaVOR67ewuc191R8sI6/NAxNdpAEJaTeu7h5KnIrZd/m+3riurdNQJVNOLGvMeo0Pb9WB
qeIV2M/ND62dq4ViBEN3viBv+1MBsNf0IJipuVJZaqNgVOoZTWQ6POE0i2X80PJoVMDKMo3HYweV
XU5yVVWybB6K7g/hKBgLWQexkrBhsNvjiUBfWhT8KFqRUSskm0vPW1gTA5C5+WFmECU7wUBPESdX
pzHHWI717wKe+5SnDfGmE36g4+XFAybF0L+1UsFlCTfwjKC53zZ59q3+BLaPSn/sT/ILOnFi2M46
MsZzA+3fYHz5mtafUPLiKFtYHiWqJIM6QXxYSgAlT7dPYoCfuvHYxVIHEr9h5Eo2Lv1lY3LyXkBr
noMGpLwcu9rdz2X7pYulO3an6njA7kullY2GkjTxJ66a/6T3gU6f9XgxRGVPq74F43TpG4FokBHJ
C5zeZEOIrWtPD+KbG/JmsW44hDYiiZ1b3ooAEwiPBRddG5nvLPVXQkemtb5Zevseix++Mixip0+9
HZpBqDvxkUWy1xDs0oEahLFUWKCKWnaYU8b4fzMx5j+vFVuX8LQW/TFgpDhM7dIcByr7En+JXMnO
mJy8f6rpCj2GLEaR4C3H9fMYwcbOtm4tOhPYljGf+XW0cWnyYGxvrTFNK089vL2oKbsMDGvDlxHv
/cADwXwCHccYkZ7EpnpZlXokLUQkHIXlcjbt/5YS4lpEH2+Fe5MdqklrZck3C/+Fk79mjE2vtxgG
esfTiVLTNucEPzOnWFSnRamVEV/aoeHc1ZfZ2FJobEoX2mM03L8vdhupSDg90+5+MIkPGis7FrNn
UE3l4lfN/dGodmX637CuFL1FeSf8d9P/SnyucFD1/m3SP5OU/4LzxFGaBWhz3bsulCXYEZWALBpB
oKVr1VtCPbRlin4WU9R5eICHtsZuNLh1Lgs9XwqgQafeUNKbo3lxvFQX9Thoe0cN7XYh5dgRJVob
aQsQohAe0oNuWSG4sWKsSG1ryI1ZP1vIX7oRzgdvmyZkaMkkmQSfvmiENuYzx+CH3dyKI6Sn90Bf
crSOR26XA2CaDv00NZLudJKyuon/T/94J39Ed7qUVOHGasyxadTv5Q0ehDUu/i77/MPuRH4dyCa8
GkcbJK7fRZwrktndaVE+/ySP0SOZrQVVMXOt1ccRNobrvdCQxevNNcqIqn7JZ8AAONg7P1riOn/6
u8zl+9FZivsCzubqrRK2ZbSmYfXAkvbbaKw2O+LPzk9CGZBfH82sv1jv8xwh0Sd6zU4og8zyqXQ0
Wbr+erpujxQ2t0lf6o4V8mUKCTs4qT6LVB+RkMc4W7l9plobvMTVdrAem+FWqe3MFMdDiNJv+7pb
VTBUFzbUTw3SoEhtaxXKPVyONFqCM3rjbO5ZlduTM2SKGklIEPYJ3uAMB9fbFXElAZju3VcUwwmj
VzMfZ+UmqiBU1zrbaSVcXk6FGmvO8+KA3yCvWGVyum9lvKQsggT3+DbItCFfaQa7ox8IY7knT8ay
K2ySUjUJIFI5ckG7uwrV8E99YVgeBatE3KNao+mNhqEj3dk2E7pUihzVk6eeO+6BHMmQX1qe1iNc
yUY3fTBAZWWEZrT4NJanuhIy0kzVigQhWqkQuvEPMijmMZyGbmv1+KoORyc0mlSnRlCTpu1+T+vk
MHPiCmKYZVwJqvgM4P7mwwIj4M7KzdQqwmqVv1osY/QqaezsdAn+Ow0sHOqMuenKGVe2U1UXj8uS
hxK+MS+jXEzjn1Dyc+1kdspKFS4X22NSijY0d4zmV1K+7eTQxFtVjVyRMaVD/62JYQdCN9xdGeVf
r4GH0AGLrpRkvbC+M0ccD+muFoaUQsWtd1WdnhAcvKWhl1QbW9ADUfTBOK8ydRkpCOBGWlkPJxxg
+/QQ7xL2uNcd9rIRWcsmZm1/KBZX4AOAYPGO1lx29K7QJ6ksS+E/Faud7AAeqqvoG0mDZwglNVhI
TaVKSE/kf9GMpZimDV8VrEaJwJDn9tBVjgCN2VstC8WhK8cJdXK3PGL3fhszR32VS/c0l7IH9rgN
oaYVtBvkkBybAL/7U5Byw6+WEft+VK27GfEVcmdkoI0vMf62uVIrVZ/DEnW7elH/Jiwmlth0wkq6
kaJ/mXUTH9/ijC8jYWSsUagu6xVVRGpfWnWXeylA5NjJJqfl60nhV+yTQYKw5sOFsn8Nv6Wz1Dtf
78loNOQLnjUkjaplSrP5UBtDdsMeAyqsoRI94BYs1elQ7zF/Q0kLACuIWJtgel+NQRcqPhQ6nRjp
mPACABxoxS8lqctVDAeGMb1YOWfE+dLXm7VfcQQHOa7NAbzlMuUhxV6dV7RLo4tdZxCFZWBM5lun
OUsIDgGWjI20FKyznvSoBIGGt7G1WkdvkpopNbK79lySPIIp0coWYWinA4RDtjQyrQYSLb2wwtH+
NUaP5aadpzaRXUapFCzo8j2YV8PK/dUO9xxxSX8VU4RDSmsa6a8Ih5P/xpwOEv71Sm4HTms2yOjI
hxjTYYmbsrz/K7oVO9Jr/zL60+jAXtY3Cv03bvX8OM56A4yu2kJNSGBcXAifdTpqug/bDezAwL+A
mBKZGdtdjzTWmOlNE8yUqxeBRTCGFOidRx+C3yfDPS2PsUcaM+DpqIPUerTE/CqY76rXZY7qEZBd
N5lsy7R7vmyxRNhQE1/f9iIYZnHkVg3i6hmf+CDUM/0MGEXLFoH75eUCkFlAOphxJFmQXYTG/+01
PyHyax0gxHPE/WWJva5Vpa/5GVjWSN90nfyJV6whAPx9C5gm362Ier3vGMFxgvRTW7m6tmH8NSLy
oZNs/aAYFG0BQ9wpn0oiGRuNIX5Crwcy6JVXTqUC0cxb/bXeJvm4KDzT74G0utjZ62LHhtfpbj5L
Xbz/lK4W+uzkbjA4z67se2xZGNJsaCwq7V+YmgLlFYi8q3cMgV0trYyVNJ6Aew77HDmYnfU6h71w
e5S8e0ISURkg/CLWidw/PirOVBnjM9YTKyt5Al1M3jPd3xrC0ieG3oCCr7G+uMmJIP3hs0pgBJtv
p5fjRTCd8HE5uv9tpFS/y/ro4hWJB4zGSFKJkyZi53QiZ+r6X2ty6vrWdJdGD/b/fcmpy/cG42dX
0D6XMh16JjOkGcish3fPXBVcQKP9Ue1VupOCqLtzVYFnUJX5dvwjqsLhU+VmKUgGJEGfubKxtgGO
XF8IfQK4FY5RAmBXX2fv6SIgK81nMStLWLWJ+6flVw0AvGsAGZ1s0t1y+j8O+rfZxZ+iJfU/j//4
6sc/Sr0ourhYtaEpppanbdnApyUCPEFD/9Ks0gWhJ2T5kf2pteSeI4kWZ16nGu+qhRDyqm+a7BbN
cvXoX+p67gkiCsZajPXrLSYKOj2BsvjDRhrqFaUaaIPITyh6wp+XyDPnEqJAAvJhzMgN1hk5NEGW
n8BOu7jU7cDcoxUGLlkwrp6jPH/y+Q9YN4TRpTk3NbAz2rNs48H9TMpOUYvny3mDsPHTgMDBoqds
yJp5QljG7A28e2s00csgb0QII3mwIiGurj0s1ggdZ/uwajVdAta1TWwWpkJ5Jp17dRVXFLB3uAjZ
/dJs3HEmjC1KYa7KSCXnjr82wqprrzlkeyuhJ9kr2QG6EKU2s9ZnXXnoBDF0pFGHzWLgRHOoQJm8
0tcYVIvE9Jo2TUVrpG6tcXkWIVcCSUzPx1P8rqiCG/5ChJ5FRRbL5Csc4MHyYh/F/6gD20lDVUtA
N9jLUanM7ytAJLzKsMpmX+yxnEAcFYfv4crmvav6m4zQyOVcc1lPGSpb8Ili3efzeJnJw0uADWzu
SVtPsoMwzNyfUryIM3JWV7efck8cOLIVbtqP9xhyxEe9V+Jmrvz7XNFA/eArl+qPhmJpzp2lsB3J
zRn9HDqzFEv63vfO2Nu9wfyckTEwlmccrcBH2+rlf9Pjry7w+SzSqME4Bih3MLmcNSia5ncbnbyB
b8EV3oU9Bv30duIhsRG4iWutGoEWcUEV0pwPQjeR6pF1Zqa6JvYhQCv8tdPa3oCHSWG79Xlv7jf1
oXmXROhErFRPDB9Bo1XK2OcTzGkQ8k7F42ptd+fDKIvC9F1vJ3BX5qBC9cem7js/C0VqobD4MC/e
67c3eHsK0KTErQx6riAHxHTSJZxvg6FmuLoAuUTO5m/yABTArTPGLiK8zWwIorc0FwW0PfwadnLl
nHYVd+YHQHt022RsyW1xXw25HsK8AJ2HI/Yv5/1CAWf/4artXhk4ps8xWCsqYIP1tf7xXpSYUVqP
WLsuSd4/atSFavyUSDVeNW8n4z2Vop8RfVGfsn2CXYHkH3HJJ/F8CN6Bz8I64pCyxqqpW5XXX0i0
CoY7zoKGVGcVL38npVNoz51blwm8nG7KPIeyT+z+cPd32ag3P3ZLhUiCVg/UZbK0qE63i4Es0xqI
D9rvjLiq1w1L1u4rR0eL7V4blVpa0PnT6X26XGd7H3bTXULXANZ86dR24vQ94pxIo+mk/IYgQPv6
RaA4YAFKsOxNH8Nz9wXtEHhmsIzlWfjrMcGhBaJENsD/aSvkdXbVl/M/y0pe00grOnGODcCaSR1H
a7nKny9SdJArYMAdDjWcLje3vN+O5C6lC67p5h3ulQ+Yi3MsxA8mgu/vplWMPqVZqSjD/o8tIfJk
e9RD9f9+VHI2VA+Rr8LTWjCnKP7gwDiSf1yg59ISqQlM+dHGTMJvDLCLkv2idhBD2dIzYoJPUNh5
YhHxtSsvttKfu6iH9MoHgQpoYZIjbSt47a+hDv/Vmq1Ril/oeftxUhmxzfzLRFrlJu/Wkp6UZI5q
ZuD/o9TDYBM4gdAjdw7rrDRaYTza7ndSoEWraJGKXv7i0Uq8kl6bQiIqrnQLpiVN0FDsmFVTJE7q
KFWS0NRVrYjacQZ22x62duIprAkCg1JO0pO3oOHLfytT1DKqkKSSGu63EBGoe9wVCmcL59M4/HUR
DP+XUOso3Il6A/IB8EKnkJ9etbeZJcyebkE2SgAMT2YDdb4fAZ7iKJ7se3RBm9cgbtghg9d0+syw
hWgipdqUHSCtzlxdZgomw9egGwmWa6U+uU00JOj6HUaR0mSWD2VxjdEQUihEIa9CRjGAzvrWy2KS
wJXBZeloZr+7WBTkMHThsVbwR77z38SL8Vsw+pufuot8VAfKQhbMdEsDcLFF+ASB6R3jp49GnkD6
7aWawf5FGBO59XD+eXKCmLVgvNIfvYQC+IEFUqVHh1/WQnc36x391PZl77NZs9aMxS8qEOKv9kGu
liqPbcWOZaZREd3l1mHKQJ5Kiy/O9jSCismNz67bemzjB1GnY8VG28p1D0dA2Nh8vckSqeHIwp1q
wJxmTzowVRa0fi5eIkJGJdTUBmB0Vzs855p88CyLS4J3AqrHU1eR3Aa2YpP6xi+DwwvYfCLWH/3h
nEIjIeg5RXWfj4evjBNdyc4JxfKXhUjotVVtaa9n/HjwgNPgfkjtoll+ajlVq6rd2zPuJBNlYKVv
XY1bR65ppIvmmIZ6UViqXAqABvitvEFijzZ6wpYhvywQLJVKdUPDI24oc/vhriCdRI36DuNY/jWo
XXPvz0pmljnskKC6B+LS4zbjrzRC3HeTzVkQSrnUWCE1yalHRIbPf2Q20fuMwuk04CcrNRcdytP0
JZJxuwjT4S4v5os+P81QXUsmyR5R6B5j/awzPLzf+Xww9MURcFmDJyDrsepxXxRNg84rhPz1Hxl+
2yCa/KDHmGVNqPj35WGmsgml+UhuUZ+GEPxqedPyK1VzDAbMctgvK9QcjIPNOaGvGl2iCFNSu/oG
PQsFCz/49a/V7Hb6zQlNEBbHmy8c7q1tal3CgyxJy4scShm6ZTzE0bzU8CXrANa0Nx3jNWIjMQta
3kJd5wTuzWU+VlISoqoEEhIBJ8DpWTU5Nn5wggt8CWyNCKiePRE9tPuxhHbt1TGzNqoqCIyPz0Ve
UwjJLL9QpPmWo84Q+hlcZwu04USsS6+BmQk/ZrBetslB0CjEKgh50dkB4QQ0bJ/LncDPwK9jkvl8
wYOVT2+1+IFAZyZHMAVdfuJ6b4M+Tev2K408jSE1/uiUztdB7gYf/zsdisVJaXcDqhDFd70JZGKi
ktmmmQVCooqu2GDNc1tWLPII6hfMzT/JvKciAjqKXJqBiPkr4c6flUlvyNITBeqqiw5l2rgwCc5g
aVOTIEyL8Zif6QeJrSXoZKuOvk04ZZbX0wqkUVDTuUhdt6ncHI2T19A9O9AGRp1kOXK+nusXq6VN
s+g66ednE4XMvtQV3jIC86mddNLywwIVkFNnnFF3BRkMXn8RgGZFdybjvUEPMRvmlN6ZZHuMi52b
trgMfiQSyIzNNsCKNdt1E8S/TxXxw19PtFg6ezPmlT5i/TJZTtlkMELemBA3YibBWiMIG5QPn/mJ
DQCE8aCFzdJyi7RLE4yN4hW8kYJBVIU80hRlzk2vtFApkvimXIeolssc/Cn7LeraJDgvoaSKK5XB
2NqWMoik21hfkE/mCPqV3WJiAr0ETHEdz45kkTQty7Y/Wjtmw7RmMPck5pvBoQWjVljvs2+GqBml
dQ2yM2cALJv+CPraDwHV5c655koHO/jZD/jWVEBAj/8+9ZjiG7FZ2JK++ofMim2ZYFAd+XPAH4me
/5PvK0cWVW7udL/f5vI/qRe3lok8vzgXhSI0BYEfzOQebcsz3NdIdgpp6gMN30DvMOLtyomnPRVl
to9W2T1R+0K3XwwNRYxFR6oYDMblTccEJ7R9V5Gez4ZZzhYMpbh5kPqtTeVoJZRl/Wq/TtS+H2rg
qDh0CPZHZS8yCapFBIyVRAXEwbGSV0RXqIDElooTLiOgwgkzLMaDFk0q3ce2U9N8HVHf5TaQipFw
hEWYH6sUlU+9RLbKDw1e4amc3pTN9l+XPhM28hhdBrkqx6mhiIWL7hCuB+ms5D7TUyMs14TG3iXE
QwmXvG4r7yXrVHUK6uY5NykVn3esCV3MsZzbixd7LOY8MhC78BgKAz9mnem8ADVL8O0iRtFOvH6t
VCh2vW1eK3o+1zcoeeTxe5/4XXrvRJZ7zKr7+OPd4UK/6Lf38z+w8x8w+TivQR1D6dhCqlRjz2M5
hLaWsxETql2suOCoiQOomgRqps7kT5ycoShpOAshQ/f7Z7NoXFnQHHloQm4eJLIhe11cPUAvn+/W
i9E4rqpKX1biTumPF2KcnboqGBK/+J6VTDjzvnqIOj3SQOWD8ZiwGrL3nn0BuHoofVkeB0lsAL1F
uoK/YMyDSZrwIMeO+nVmCOKPT5+m4PQsK5KMBmnh60vhIO5jjIyU4dbvHEykDXU7+TCzB2rEyjyW
dIsBUKC99skk4VGuk73GHezVHnVymF5k9Z+QDKgKlsiMtlC0uejPq23GWtpvADc4H52NhV8Rtj1G
HXNXQkdXhQuQjjMJHZ/vbWYrEZ3993t/nNOcJvw/DU61o7yvNdwQRAj/KBPb0/jQZo9xb1QTas2g
Bkui+IgcbQg9pF2aLsDFN3M7rmg8sIttKpivFbvT4WHxg8pnEUoUzn5XW5bUPHy9PD9pw0Horb4v
KUeckAhiiWiWr2rH/HFfZ1RpeRMJajbhQRnRoXsuWpzRdCr8lcYs3VtHrnqMbPH1DN9r5ak17GQp
If6/HdKK8dClfXD0Iad/SEgJxImfKiYJ6w4VzvHS5NBBEulf/XyV912EpUb0cZxYnNaSm49O0EhS
nR6vW852iiWtxYm351m731TF1TgHJ9nHUZz7uzRigLZZP7RZqnNOsc7Sdwj2i0ASzcp/dLhhhWcQ
mlgadq750FAf20jvqogKKk9TPFpn3AZ+VBpuqRxRTt3Vvgd4Xdm0dBYqaCEUQMIPJ2Ief6ufLT5C
okOIKOVyuiThHS2WSn7/QmUDoOW5HrBelj2YoiotsoWn1qsRreyi1TkbDpsz9OeQud+3/Re9gtkP
AlDw/e0KJGuVvSHweSIN7LuoFXoprTXolh7EynApmqvyKtsN1OvEYDI8bsJ7ZgwBZrsk0jfjpegX
2SBGGLVlD7AigslqC4C2doLzrcGJkzVOg3aordkqc4bykY1F8SmAtnWgUgu87jwFyqc/Kl9bALvj
hHTnjdnXozOemAj3X7/Je8IaelmIZdiZw6tvVjaD2VFYjE7VOmXnjaxpNFLLgm65CfDw2n/oxRhQ
TML0QmN3HOZbx8ccFAeM84jF95oBibj98/zv161Kn0rBqZ183QCK1WlSY0F/zoowRi8zMXYnvOUk
pL+rGA9pN07Wzwd3OYUaQGS0Xv7aZRs0WWBqP31ihjE4h6ZyABjO2AP93NazYU6ulbKHO7qMj/mT
rutoW3Xj+00l+Royp0yZrNQB93vymd3Nh4uQrkn6HjjaNDMWOYGgibMgKLkkxPvuSHirzlV9CJ1s
Wlw8eqWTNLSUmTBBAPypzd/BzIOVRm3Wq5E9piNFrfHh/f7lX0NBPaD21+DckPpRKj+ZcDiSt7nB
dnPG4QAeOnR2MgUdt1qGNnv5Msv2NIvEj1LYxovSZ9MA6aW87m5ajDIDdVxfH9B39rYsytnoZM4a
iTWV7X3a+X38vOJvKXuDwoHsUfsl3u5zzW/204p2Tklhkfvg4wHF03deVPe6Z3I0LuqDxugck+uw
KiH08K/3LjyxD+Q8sih2IaFCnFu1drsXe03H3gBGw47ZipgQHkju5Om4OTCfvqqCQAdkEmPFlhYw
yCxYbc8WgUYYN1d8kLJLqRNUQ3q2M34UC6FN86mLi7rhgBHA4yR5SUPeQYlwwoF6hBLBmKIGQ6Z0
Kad2pN1gleVUniD+wfkK7CKn6Z4Le8kH2Fuf5qf3i1kTmt6Mtd5tGVNDoLlc+Bv8zxir/dZfpyec
eCtOPdcvvFJdrr9b7t8ZP0swZoaUouGBTnwaW8vJczvaMvcjKDe+56bEZcSMnXXkEGP8z0NS4ZAm
XKmjRgvLrFlTOSp47CPt/m4cXS5V25VGYxTMAGFw1FITjQdQLQZOMG7Yl3NgC3OE+CqZ5TVs5H3a
O6Ri7NDGugydZBDYX/18UC28LQuE4rtlPU59CBG9i+2DahXgVGDZJIeSmYrjcD2qBysvX4jH1KWn
5KEgr55l9ohi9Ou6YkZ3Hb2MAec7trZe5aXp/C464hmBU4zkV4ALbM+vM5ed4LvxrzZPqoNdlYDR
XH0/63mpwVaME+IKnPOUmSIXVnsor6O0+C8ysY6GRwLz8ZN0e01Wi8gEiPTI4RLqsvgQGYHsTDK2
ryRk3iIkIiU0mlKFM5mMRNeoAMCEUFzSGPk86EUnJs17ufjOaDfrUUcNm8Q/zC+zB59yxCwWliRW
HNdKzY22BMeISFyEY2BMpAvmpEX7ja2IpjFPMC2/E7C5eVBbHOFua8jMMz9r6QqM5tzhXPhiT/K1
V8gcOz87vyDXjpCtIafU0yScZiLGfy/JSeo9yfyFaOLGsM4zNRQeNkMfrwh2BLD9AHk73P7aIRkY
fSL3c85f1n7AbpJrEotKCIo8fevbtPQjSVTEDFkvZRaJidmuK6iD6V/FSSkPwm6jqiBD+akBQ52g
o6o8J9Rd/PPXZNifEFhBLKd19mP+GNy4so2d8qA64iYe+rJLbVEKXe5wctd3c2EnJcnYvRhrJsD6
YIAMe822dFCQJbtdk/ZjsUfFxOVxNv+Xnea2ecqM+VvgI4ySMOizgoZqdB03o+hbf2f7Qfd5KT3v
e6pFPEB9Dcprvqx73lpu1NBDPbW2Q7sSDZYvNnaCzLr2nxWylH6qkG8/a5EALH7IzvDjq/QISwrI
BpRu6q/RdosB7KYfir8jOtAndr055qa/6DdZp2k7mHx9UXpSYdx0apfMWC8Sk9MhqJ9oaQIGbf02
Q0s2FoOlwPtokN3TDzNr8xOr+HSlNMfy3zyxXlOt+PDZ/RNAobcd+dE7t3rmW9qsEzexgY+dKE8v
9oVNkzpUkjmze861Dm8csg4tYo8zoxwq/Pq8K3wkYLwITkBiQPBIvqmFDnI+QUMZqIaWrO/p2E0a
uJO0QAnmYkKMazCtDA7cdCEW28Ost8xjkY9WZmWLuGsyRca2qXJBXQYXCEOwsJT+KAV3raa6m2VT
ejj+j79S9NIoAD3AYcluVyQ6Rf5fIfN0anhN1njwx/bHo4zSqbqg6Sbo+STjConcLqKV3wwa0Xqf
GY9sFOPxVz7uKrqXmEqhdVlD1MHMRFUiH8bb4dpzU6jDFc677xYyia2wjpyb5qIpB+VnU1YD9nhv
8p22dq43c5oDjZ5oDGmaWuSrwtO5k/NJX3IBM8RtNThJ69pehi2GCaeOAQdNKhnuYRdlPBG+D1zB
Z2jzWcSeiZ3gAkt3Ss9qpHKmno+Acbwtj+AnISUE/RyL/l8sRV/EAF0D420SvuQGXsCOMIyuBxr8
HiQKSSoVFPQVbkdHhVsqRxrbMbPojsPRKprBVrbGppFt0R9FaXWvW9YSEUIIoyF35AQCKrHbDlrw
KAYOcJmVjTJO26fJ3WxpKGJtJrEOjCQAppYneZvJQW2WHMxZup0PWP9MLJ6SSkto0uO66WbQaUR+
PgyonGZBFSJnVpp0ahh+FvOQiphEG2WyDIfMU0yMkRM59DrpJDbGqM3mh7UP4BxYydN3AMJhtcJe
avu78IncgPlUemY9+IHLMzgRYSYVEZDoI91HJpJ8HWk5y2fwXwLCQrjajr1OkNyqaDd7tG3ga4A3
TywXZ8fg7iZzlkWi4duhHwgzgfk8agt+N9i2EADBCLcIPbt1pETpUyF3ejklcrKPHmUuKNLw2CiD
MOM/DgLnRaSBYZpZkKCxJCNgYMxsTmMka2wj1f8IGGTh3XLPpGbktL9quxjO+t8OFUXPPjTGnxyr
Ux1Ad5pwcTMU7w9zITd+RuYbqoXfNrgNOQ80QIlQfDz9bJtXVABYkYNsJHvq0hj1hEY7DOsT1QFz
ArbcBQKQJ+IX/c2OVJUEDek6ljqmOsUmoAWB0kzenNpRZxgIvE8/Hwx0rPi4bcZQZ5mbWL2Di1oh
IWjl1po9C10vgO9dcx15rEALyD9SaWJ2u7vQ2U6AwlZ+ZXzTWLa2ResGkW5cXemUKaCmQF7l63Io
GB54OegzJRKJ4QF2OjkubT3MidHN+BhSGYQI/kKuK71OIQizTmh2zQ8BE8cH965q/hVAKIouRN/H
sW02luR2y14hhHSQJfAz/GWI78J8gWyA/TPD4e7qfjHdKcwfnk1K3sTJX1GwBf7co1n0DV0ymUMx
62D/gmFIH/pOCSzIUFT5U/NkrNu+OyUxXBGO8ykfm4wRICK1yAhvfAA6X9q3DNl3H2woJ4HgvbcH
oumFZoFY2FE5zvZX0e84z2hB70eUDCmkf+bmLnJpMXBp/uHDwkbbA7TqfxpMfIJjjZV53EtAGoyh
m1Z66IpSCw/MeQ11RK1EyNgKHNv8peqnuvhpVWLX6LcEekZAWk5nQdOwuptrrZf1jeRD5qstCaaS
QeIhJg5Ln+29O3wdH5i1ZKj23wC4GXW5eo4bGSXDei9ZBqAzWB/9VIHHEHsUJO8Utvh0S6TkyLyx
S4oYx/P+hkWNqDeIs0AoEDWbOOaitwJpkXNL3TD8NBLIGLhxzAxdv7wDYTVx9KzTwjtYE2n4lhS7
wN6s0+GiIjnSwym8/7b1i5IMMCB/sSQ+5SNkV7Z1VxaexmfxEdsTY5qnn/pDgbTlR7ifxGthQ586
Md4ZteJiBWdz4F5JtYGbM98p82cHiwGS7lV0h8pDxGJWsVMkJZD3PhaxyzfBoWiUw9eiaQsKR55j
4dI8+xZe6DtAJ2FIb7nXuss6OJyOYStBuN8jtdp5cED12IthshMtsHCWj/TzEtADDQjlVWKbQ1yF
XzkETBHJT7GUqgq0E0LrvCBvRbK7gX0rJsbLBOGmuIx691n16W7Pad2vMdfi9TNTCGusaijK7oJ5
sQ8yUEYQT2NwGmNsepbQMT24KA0OwEFxROlwDDEc03BUUehZsp4DzVXnanzECfov2TBHUV/nmqu/
OdpL5WXxCQ2+LW4jyyV9hXXK8DekBQwsIAV9x3SiPdCzHeHfRply9meO1RzUOArJztGFAFR0fJV5
0wRlgaf0nBA4LYvbpmXofvY3fO2PTwxLzU/liw5fGy+tz55ccM4W2lAEMPEnK+oCdajk/2P2SBAa
fAY48NbS0lDIxAsmbJwrGXNtsM4rhffTIDtVYz+Bkoxc16p6y6lL952vWwLw6GOFj1vOY2IIk5Bg
D3h4BIMpO17D2k/scrmhbLMJ0UVvxAhNoJb2NPbfKZJtjXWEYeXpxPiAcgAM09UAMXEs/kGo64Dx
xrpwebWFCodVP9eQa03wQ3dtt765DDte/HU67uqjLsVwR/VDiUV6thUPgEyFYEV6+7Gcw7YlvgWD
zCbccSJkYc6TYJkYWy7HAqJ2/SmcE41Ix+tIdikIN9/wVpgGX1V1VkGdoXsrieBhtRKIb3UzT8BR
w84AvtKtjnxt8k1hTIT781efSOLc8ETXottEDMyKaLwfG95UxikFJX+SqrsbPFB/7GN9ir2JlAGr
SuDbdTUpu3GOdfbMRyIkrIjkuOBiuK0WHIemPulNMeg1PLtea2yl31Jd+14Cnz4izO0pTVSSGvHZ
CENT3sKj49Ve34SDYwrU43x6hpVleJejH+MW2d24cqaVAGxkdlK1m2/yYl9jQRP7/31vU8dxs3O6
y25qIsJv0ybAnQ1LCrpb1pkUKLl/ePc/QXU2OhUpPOSZZedT3z991H1YmRrdMOnxENtxt/QsMwKX
hx33TQuBvShrxynF+OeJL3F6sBAsX0qhfj/ioblAAfGubSQT4WboXKd/BbU8iwFYOigGT3zjH83d
eN2gJs96Q/Rxto9WEJ8/vcS5fhVbZvb8+yWnjJhTiAP0z7gMjExtlYnhSILaN2M8/8ltTN2FgsAf
gW100OVID+TAUNoidGfT6UmLxNKHikbCX7MU3jB15cDq2R5KKdV3B7XsWvVLIX3K+inDbIsxFcXo
jeyQ/8NLzbMVZMhv1ZO2tVpN3t9+jqweSSZmgd6E0AXzTgtq4nZ72MHwTS+F5KdW1rSH8SeJxnKh
PEqMGlHnw32gK907bxDrxZC6BgHOS9JvzLqKzXFM2OGT7t2TJ2Uzmtrexgi3NR4NtMAbAzcMQURF
UsbGC4pqLBeKQL7gAgNrdRrq3VkL0frb4Yo5Z8T93gMmpwCYGK9oZzo7nuRquLRw/cpR3k/2HE+Z
BCBaTM0PzQj6n3WBT1QJCbo+kSyk82B5DuYto6n1n3r0vSbJA/J30iU0OKoMbu5aoAwE9Z5KfR4Z
5y1XJyTXp1DzQN7u/6ln7ijWEgMt1LWHhGPXmCAuaNI9SGCnmP3MRkKlCzqUPuDBP4SXxJxSEXbK
PO24e/vMfcrWQv6H7f0mEiDqnrBqo2wPGgoezeHInJZd79IKw0yMOKM7a8xCira0p73ROB5piWsu
bJJxzu/1TpvDpxiCrhGPTTF2F5HTCjZf7K8L3XBxFd6nDLqkBCatfAlCUF9Rf8VYeyMv/fe7zBHE
KQdzo+fWKrZ1b3tEjhBE36ap6TVKW7oBfwGLM/jdKQD7lC5A/Jmq1YbQ2mn0cpofC1/1O521+7Al
E/kDpIQUTN/D3eTMsJjct01Z6Rd/+pdKiBg2CFJCX2EuqwUCOu6cKpuP+dDhqL8jj62mgZAFbfa+
9TUhqihsJNA559P/KG0DJffB7o0ZZtZdCXjCCq3iC8EeRBiG4l5HbtAeweDPrSwIVl9OhXtOtTAO
ebRFiT3RU02Fct1cgbXjLFq+2gN8Wbr75A6u8G1Qxh+1buGT43Yh+U+w8rflGez9L1eV6ysbzPK/
mhw7qrMgp8MJlpmp53BNiSmyzOPJSSByjrderxFd6X2jTwgN9z9JxJV7mup+5rtRPUSS7esiQK/Y
/o4GGIR+cP5RpWIqUQlLDsR7cJ2xgacMjAYjRDjkZWV7P59qH/3dOyux+Mwcuj6djej+oECxOkKA
8E2D5G6wMhnJCVoMGfQ+zL1/HgnHg+fypkAuuWzg1AYbxEww/wObcUgNWvgY2V35V30Wix9xOHtW
7uovWDn5pixt3zW7FfdMSeshXrw9v9fiWENlvEpht+NJP15VzgaTsAOJwJFqMyt6/Wb1Fe7YdsHu
jip0VVOWLzS+mOgTq6GkffT/KTssFWc+Nt7olAOM/T3pJYp5lZHh6hHgcH/tHtYYvhGWMS4hmU7Q
Uyn9om8EgCvBCMp51hUhlDg90YWXSSy3zhseb2+bo8Cv+AJ43vk7JBDyxVFVtO2W79jQ+9Vl+2Ec
B+GBRTkYy3Sqcb+pgvBoMMMub6h27SDpyGPdkGnlaoVaGT8Jsp8JK87Fkx37X5jaU7OoqRwipSbi
Hga9DF2LRcpNNw41RojO3EEuQ2G1MQfKpbsx5abkX8X1aTjy28wVFAURND5fZKe8OQBNs6X4woup
3zj6FRpPCmNgVN5sdzoLLLwPafxLF3BR9eo82BIva9B3onvPNFxeLQIwwopa48v23foiRUvwQpat
rKGAWP2u+sMRqBm9sPTgKl1m2UfHy4Vb+mVPr8RO2ng5ep6paxavul2nZBOE5PrYMRgPA9h0Lf8T
dfDijxHdh3W4jGYHp3xzmwjVUTfFIs3KEqkkv83Lbua8fLgSAsxkia8zupzj042WxFkjsA10yLSZ
J97njtpohQjS3YgtFGzPindoDhpd0di+2RevjxCw61kqQq3tcufwOfTeiIGwJ6GQqwEVWvuy7H1G
BONM8swZ/xoHYhyvqG1NE7m39BMKeIqHKN1ZlTQjyhZB+4RQ/25D1BlqdI4VrzBooagaXkBmuQpn
HyZ45oQJ16ccwHCstzRRQLhwaU1cBNiRQV2FLea7kDgRu9g/m5D1Kq9qyR+a1DcivzMjyXUABm0Y
TECaGUqchEPFSj5Uu6etAEyuPbaX641rDBB2ooUrZmT5zDkKfPNGr8bi2i4jBpj67O8HL+DJMUhV
vTtF2ERowqeZIwmW3EmKxpUe2s3EW/WWbaA3+3VmghzFEcqEe6sg4ls4ATPWyqjbgzGsuF4hSZV7
/cygrJFTcwykVWHTf/PCkQG/KJhjSThge6tyKg8PQr+B2D4+bd60ifcF+klCah7J9NJd8ecJSyuB
pvjfmilGGX5jzpsU4jDxBnXeLuf4mQXYSK9s1nf12eE22w5dw0sRtSL6rhanh3HbnV9QOBEiMM6d
Zzrts6NcpyLU+pZd6SJA4Eyb0RY7MgK8/SL2Rw6KvATcQoDwhl2lXK8Fd2dPCrYWOpCQeojd8g8U
v743f2eBUE2S1sxjPn4vRaABWoA8p1TeJwUgYi2krXAasfJcRW133beJkTVmGRIXJFteSTAzwrsf
ZF1CU2MP1Kd0ivFzh0xuPjS4En/SDKZIxZC2/BReglR3p6Ic4PS9QOd1pvgWllNsWm37mC8abumz
f/Onxld1mYhntVb6NYufrQKYq9Ov5LIuSt0YBrgmv+0qAo5LiJTcjFFc2IW774pbaUH428uSXaq8
4fbHB38KJJWQSVqCsw29tJlM6qxKezOrPkeZsD0ghOkWliU30TjdjomyK3RpiWTQvptJ8bPW3Mpm
7UxN9Mshy62aaGDZ5tElo0yc+CFCz7GO+S7tLQYv9vtftwEFW8PcHLbJ06J+BASLhngrW8FjNA4v
VmOlI5B5HVRTly27RGuLALrd5xRyq5ecR/7DP6Jd0aMrtuNx5kREvZKPapoQCI8Uj+jRLTsR3rO2
8HiU0OPT4guxz44MJhpzEnTZ3w+LZYlDEGzPN+H97dhdPTlNEjvGWjknyopE6U4TokMjl5+VWdYU
5RkUU7Ivnq6haqkIoD7jKO3odIf+ulnSg4nglMUhJD1/p3ivnAVLB1CHvFO6XyZr1SVJYQ7ni5zD
z/sypWdIpirmBq2yDEllzEp1mLRWcg9AB9aTgkaapLZ1/r9nn7uf1HrnmRlpFdmpFxTeUqpiLfu/
UXpQgmMcXv1mhk1VUaak05pc0ItOcKSkXn+bdPwxGBXMgfPT91I4oH1t2KOIhXIbiM0jLCWdjQZE
8xVG5RUuYqaPufCzrsMzfdFvTbxQvpCdjkBO1oL5sZtkLUx+G7F5D4blPjGHYwRPiJiEMHB+7VzJ
jVtfXUGCzBcSk0K9dxYuKrcaUdZdLptKu4YUr3krBdXMwcMDZixRZ/aOGXH4M3o0+zgbTlFZeK6l
Kx9Tg5ERKtGwaVMCXLfrcJ+UfLos5LvCLW5EII4H+VMwWB3sv/gBQOjeHDcuk1nbKXUpvyzmKgnf
1uLMz9ng0N3XCy1q7E5OYa0UbRDdganDxzp9wtGmbrUfZAXvkuanC0IgxcwTj8awtvgyxnwWBrZg
wwAPAwsbd+K/J7UFcDwMs3r3dsMgUoP3n5SLOXqu4iivGDB7Hk098ATYNB3S+6amLHH95Poz2HY8
AEL00b3GA/wbkQjlKW1DFOrO+ifBoxIfwF7q+cLiP4wgkTIdgna/O+Z5ItTGmXmvSuCQM5YwPenz
Sjg6Lh0O1xiWG42AVH5ub4YFM5igfnVqumtQSlnXtnbx0bnYSAhTM68sJehegkuUwDr7UH58IwVo
P0U9PV/lfnuPVpgXW/SNuVIeqQRThXCRIHwzfLZ1h3gYfvUXoBX/BSy86jPndgKbPUkqih09+LJK
T2637Xth5+i6VNJ9HOjWo+o91QbivloNxI3rbPYV+dB/thTGdBNDgt+u8d8fVEWSrvd40pyDIFQU
bs40cyb0h6q4vFYfAckJe2M7ksXt4Xt/fturf6pRZvSMCTeKZfb/JJ0w0JJ8KdwrDEWscXBOK1Pt
HOH8Z19UsAb2inDfDdFzPkCb/rOCXkda4rUTu1Ekugbe9E+vR/brpNYZrrcL5l+z9qdDOHUnTUYJ
5TieIwS3JmUdwFtP6d3cIWYYX6I3PUQPyCpZE7DdIKlQ2+6Crni0xhYxkhj2V+zzxX5AozZ/usa1
bKQ4k0+pbIPZDow0yRia711AbhvE6e7V3ywFXjK//sSZFM8tpTnqU0kqvudeGAB/V3IQBpmM0KIa
zT1ooECn64wiuuCI6Bfo8BMAAitrgyxVsQlp3SfHVkA3Xc8t/tU8RCDcox5tIItuF98B766Umzsu
pl0f3zdNeloZPM/6ZNxbARu2XPxGcfqcytkcHtZMJEQgsLZXCkfKRkz6aJ55WriXTJlZ2+OpJ2RW
eBa0KzYipHJOyTiGnWm0REmKZpWAzWvEKLl3QfkyyUVqIKiUGS9EM2s5jJF49z+kODfPT79aiY7N
qh55YT/arLO0qKIx4CWkoHPE4+NcMjGRpZNI3A4gsj0UAsQWA+dR7K4JTAgXcD57BmfejMj/pNLc
QxDJjdOI8WdPRLTjltYWc5+6YZzPmwgrchcIQ17vTFD9b7PK70m4Dz/pUYnkXtafZSgf2EWpajEs
6lwHcChOj2oom6dDIEYTFL0+jQxjg2hFafcD0BmatzYcJnFyxFyrs0XXrNDPqBiMWLb8cI3zrCOH
5JMgok4/oDhLfBK+HKHNZj+50cclRHbT3dAYHYxS5rCkfYpWxmME537PwMhlJ/oP1ltlc+cp1HjQ
nR647FKHyPhbAJkWrGmTtCQlaCuz/kO0kFcgxOPu1RR6n0x1isJuaAXCkhwELJtT2wM/iPen+0nL
yhEQ6lL7FUhMvQeFhjZ41VPOBzDR1hQOWvjkvUxJhv2N0B8UxMQOfSck4BnI/rUlw/kxo9/IQGc2
tp9h2ydtRYGSpTnFJU/ymqYkg7Yeqt+whMI1vzAVsRwBXqtfn1bXCOzSPFe+eYTyyolQ8lowV5aM
eBuG8PAF2IkITlBQYp//gJOsGE9j2NjdYJxFsFY7lIRAsHqYZQ35Fw+umCxscrEmvhPXCXAyKdJa
m5pVXnnICYl6MFRuLmFyOzlL1FDwiB6Tz3IgFKmTylT2YSqBg/gXTbdLCfKBq6IKUMMQLMj1G639
1HqLryn4ckJX6QIzWtiPUj7yxJP6wc8zzCDVQrItAgjvZUjh3FJsgaB33AjCnkQSlDMdZlL2iTso
ihdnfDGvO0IlNThFuW+/L/u4Mq4h16mD87vJKAocKcyw2TgnqRMBzBiIwNPz159B7wJCB0o0E0FQ
yKWMHsyx1ZTsbWPCN1cv+dhfwoiVtobGmu6IjqyEYXUnBiE8Ae4lshdm1GrpyMWbMyOMzXa4+qNf
pxzGzs4eYsY16B4x9TiJdS04oqDsu0TojXrLt/YLDbbxm223uhIx1rTOmq9L+xZ84pKXfmg4PuGF
uN9z0tiEoRBnooi/wCeDkLwUktsqA4IioADdBnjKEiYjzRj2B8FnZ8Lx5GnzuD8tlvIE1kxbfB+o
z+0cBce96V5uXmqLGyeYv2NhrrumbZ8LIEFcIxIGXDV/qmwKuDogSYTiqngMyZj5+8BP/x8XFSqE
CnEBrlDEacAk+2ejux+72P721TIncpm39n8op8f09k3+5KVmYLQ1fH3+3wucuFWWN/rXstb9M1Ey
U5GaTBJOToSMlPoFX6+ptp/E+23dYijw1C9ZjEOz/7tgeyJVISvlDB6Z43KhkyyvtcX9gby7T4pt
tpLcQD7JtzaxP7xQJYqTOQvBFdY5bPC0fV6ZgOvnM140h7jRHj2XR/t25VYPItyh8dqN8ortv5aW
VOGsaaYLTSPzBsWKjPbe3ciB5C7+kUy6shJwMS7X3mF6eugx8YvK2w/9KfiVi18EMnsp6XAFARnQ
qbureR+jVN5ULDivcGnNH51i51/OyPonr5Qhcw78Ii5KYGs6HZq5P8Pt9oOlabtSksmyCNauF2vt
i8VZpRtwjZzcWTPuGSvSi/GKYvawo5A61qRO4Z9gAs4sE90wbS+8zdMxbaXu535LwTv98E+LaL5+
uga8wAoDdtLmqVkVuWcImYUydnbn4a7rTcn0QBhytguppBvboE2327qZrXPc7Rsa7WdiL3Xi/N9F
JRJgSIOhvVDTjMjhLxFv0tIyaBEzR8+0VmjKrPqk+9VCwhaorH6kqkO52Xg9s8ZGoW7lSUOtb6ta
ESbyMgckkw4ayWgYc/JSbQ5f8yJ+6jng0yoNVPVJpv5azEahaSVdLWARUIW7Uqngu2FvigVxJ1xe
cvheEGnaGMEcMJe8Rvyfw8sImJfO/WAFdhDuSLOG8XsEdY3z01ziLGQAXFHTGI9lINU6ZQwhPHhA
E1ijLkYCFNBlCukeVmthceU17CrKQvY9z5h+iro6T9Pvs+5SZwx80h5oBK6+hC2qMDiMLrDLDmju
TFsbVRaPfXiEI/2p6Wr5PyTKk5DrDjfSfYwlrNh+aVwR/f0fN9MX+VT3WKOpdsIDD8W1czk6h1xg
wnm0mgfkZbJTfyzSOpQ+6YOgHctVcaOEzUbn1WriPWQQRGbE5576V5X1SfGMQz4Kzyh0x+iGYBj9
4X00d5XxCL1CXBD7XRGacRhv+dmXmVFvNLzRGfqGdn0jeJ/QRBcqysWKWG0NBjwrWrDG0iI8AKmg
QCRm/CRddrwlpQ0YJNzCuVhH2N+9LAbiHByFO2ua/4jM51nulQ5ND1C+5aqGJEXYEV9MGlRwupOc
DOSSrWNAJIzEZXHDoawwzJysrHBfW+q9uDRXIt+R0BUzSgwfI4sZIiB+4fDlMh7ItO/82AsPvm7v
Ot2jiN0aISWsfFnBNMIRP7U0B303rx+CPREDLTxlw92IB7tcWvUD/qCqMrUO5MGaSnaJR9a3deDx
OICMXAH9dEGsMiulZyfLpE7xQFvQgz7/gQiEgoP1IXxOONiAZ5fJhaqnQRuaN9Fr9JDcxz94LNNl
y1Y6yo+QDxu8VXS/aIJlytKBHpDspEO5haL9vcPRdrK7/n+akTlTWjOcr+VlP44ESQDm/ohxDQg9
Frh7CPMcqF4XcPD4Xb8qTlXKpnbxi785QRQ5rW5wz9MnxDIhrAsz1PVK3lTv7dkeXYc0oALPS35h
xo9BRzusSiGUa74374OWxRd5pgqynBsxRI1NCseZKrN6xG3PnkdUFB+8AOhpcrIl9vF3w1vPL2WZ
UR+7CDNvFkjbtVEmd9obB273whSJ0WX/6qKhiArCGpsA+CSY3tk65Tn0aFTAVYTr46KnZDepY7Gj
4ayoFDBjmcLL/O7XGiwNxV04dJFwgFm+4SsYyvyTDqbtud6oLMrDiw6mYnp0TGYDrh5VkBHXJSFe
6De9AZ4QHUWYwPkqBID/XYiLL34UrHyRTPdOmWFpYnTSeHv3rECJ6FjHeL18hi1gqbzuuOi1QmgF
EGYO+wzdhz5TgP+SoFcvxmaVN8CbPEMohyrH18zcEiGFHZcamn+WyMc0QiSKTTQUNM7SmeHBEovb
OHNkjyo96N2gpf3ydlefBnkFf4QVhvuvhXSyMeUZrpWwowTof1m6HFhRIrKEkfc+634cfRiI9e/I
WLArawJtzdGYbyODy0gE7QyA/C2uagcWOUueP/mxP0KtWTASeDdgAXKmBpd8GzOawOavULHSDWhW
oMJ7jYT/0KF6sd/0CTidH23aLTLT5OOXIWz7HdueJefImwpEQJpsm+zficIFSEcT6O+5u0KEqgn5
nTNt1x00Nz+n78Q06E+wSCEXcePweF025Pt200TvPUdbK1CaarXPNZblkDtckBQ05uNKkW8kd99M
Lccs9RGfnMpVD5+AY8rY+Wiq7oGNtH/M9uBQfa3cjgCLLqTvTWGrJ55bHzQP8jvap+iSLv/MSKta
HwKQszDtO5EQIxEIGr4MJSxBX6GnNAV9mg1asNWJVqy6B+EF1wN5kdgLayiPdPutO+AGoeRfInfr
OxJkh6RLgttneakHlz9yNZocvV5q7vCb+Gf0p55MI84ml+QvLhtB3iowiIlRpfONm+e7MjoHuXcx
2zVdqcNfWpVVf5X/gJnO+tcRrGiUN7FtgFdfPxS0VAdBpI6GXX6YWGlLS9WMpZ8b9sxr5QdzrFfb
fC0s54R3LwbLIshgsONTFU2/3i4KNIjZWEd4YJrzskVQKQ3KKgnI3CbgldBR11UC6YqsE/nHqQIb
0mj3gUZjDLWZh9i72bCLCd1AdEDLk8V+vN92UrA3F6HD8Yj7zLxtXCYjqMQORw89RoFY07VxIagv
ngpJCgCq2RaEQuj8fj9fW7/Tu/xqx276WgXm9qBn1PZe68f8OpwjrhFJZiLaZKDJ5uDQp+WEG+ni
HbRZGjv+sKy2m58bdRU1d4MfiyBt5no+TwLJUBDnlnxyynzDVkcRedmRg1g/HQW8JgCJR4AjF3Lf
N7gbfrZmm0V3HqrIGcGtMp349eq9O2Vu+TUiAP6z6oEB3JA833t2nnN1XLcTBNQ6m3sAa7KE415r
1+qu9Z44v5eNL4rqcUcRZ3tD2NalDWhPkzvYcUDGYB6te8HxWznJNf/No1a+k2tCpzNRL6Np9H/B
vO+2P6po6q8oWYpfyph0F6ChT0rBvTcIe8ElfUunN4IBFVvVhxuZkBkui5BGue4B2DAGS7JCBAkF
BYoHaKLTtYhkzlrasNSkIcJFOd+XoLHlxpkeTlTd3Y62qpDyxWRWr3zNsTwG5N6dCH8wghwPVxbr
kjwFOEFR0XMZJ7lFtzsnGr5NgfqMAgAOnC+x6nNV3+ctJirlK9cQi40KdwFwhUBQsFFE/zlp/fgM
4mvjzStGDPl6QHJqzmWg71mRiH8hpF229iVl2SfRc+6GDfF+fzCs9kwPLkX2S89sLekVGenev12s
A9PKnKwiEa05fR3BNSFzEvQpX1TzGU7Ff0TWucK3p4z9lJIW9bTznOxx6E/TC2Cs4fC2i9aLQAa0
TEWKdUzCKaffMlKOvHVHArqUZVa3+CiBWX5JomPKLU4GXa0aoxG7rIR6K9M3dtfc7/DiXNKLXbS8
JP+v1eDbKaRyXzsxXaKH9p5kC9zy9qwkoVAdl2RtEukDONdK7CjbmIgKZAatA59tQNrNEjaOHugk
LA/O9UxFFRpr1uCjGxCdPo92Wk56oggJqZMH1UWlOY39lbD9Dsc+TVC+HMr9JKImU2ScI6GWk3NC
rULARnTBAdNMkC0+XMUEZ4zE6TWaF9SU/6ScMFOsWdaJMXHH19pKzgvmIIfAc4KLYzP7UT7Dk6tP
AH6XHqBOxl5xERv01tLMSXkakoOoqkP3EHKNpRI45Pgd+9V+LfRiqGd8TSDpZiCmXQYW6kKOJwG2
ntcCuDkNDgOYIHmKIgjPfNR8pYd1h0fOn7t3Fj1+1z3zm+V0yucUpceu9hhqpNNTJcUgD7GgLRnA
G5UqVF5dIv9Q2GURChByt12lH+6HzNghGuDGKRRRN8S5pB1vm4hQ6v7a0ACOAkx+QTPTasC1nfcX
W02AAUf7lhSQPxkIh1GJR0sZwPm7wzn8Q1ytXWW7Mra8imsQGp81HN5D4GFc0zNLpxR7Abuj579p
HBs/8YKKvT3D9lRS2RJUGgBD7TiuDNIDJvabS3+mmApuXTsUIGwvVLkaXv5jXdEL7mEGgIq2b+iG
ff9nquzXGSTBg5M5jgH5iDFPDzeh4G+LkxITC6S8+xVRzv98DbwM1wPFGHDm1mDX0hb14bBZwpPA
VDR2aKg1TvD5s6EyKSCnOGl4qcRewACjiiIGqApEFZ6XNjpOVf8vNSrKT7niRWUNKlx53wCdIAIi
TxKBvgpIAUvSyD6+mcKR791o0U5Lmrv9mXATArBd5+Y1fSRJqYuBZpoBBsTOOuIQSo+UrB5u20PN
gClEc3iL1ro/+Gl1va4466IQrI/BiwMZsT4gutxYtthLBEMZlOfOPNdpPa5Nxb7y7nle2z2tQkT5
JDhHk3cbbwCq0jciV8oZoTC9bt7gTHp3MJIlqtq/eqee02uGCapq/44yfPfBTqlCKe6I23MVmmIT
vSSLM5gE4HiQNGHrcnu0FJWCSdIfcwlwMxyz1Np4pwA2D2cdQeaXCcIfW0vqcnTkABhIxiJmjltZ
VjmxXgfiFd1PX3ewZkSr4j8f0Es/T511LjYVP8HM7zdlbq++mhwkBZy4DldJnOPyYyb0+100CSKg
7NOC2w+STJudwHcvWZ2GYKyiEdUCl3oADf3ynf9a1wYRJ7SNKUKnldN3PH9214OPhvY72kNEHanw
nhch8ad+mSvRnokKM49f5Gq3S3fLc15w1E7L/+3Ms+fxxnqJeajSczuZwnscwqVL1lyf15IrRvWP
1PrZAzlW9MubbJTdbl3y0VcPXP/rTwTd4zHVFkGGdEK18VMjaYxjDu9PC4FA0bnEY+cTk/SHObiM
hS3mVprSe6u3CGGDTXlDMSfjhTRUsys63louRTLWOQ8FoYzLgWD+RbRpnoTL3j6TuLLVovFGepID
sTeck/a6iHCeGb97DIyyckS9st0e70F+zUDKYXCCc35uc6Igx3uHTwlgQt+K2WkqlJDnGXlCrjlu
nnrbDrnZFctq3X2XAXvgYDa7FIIpjizR2AuWcxUkLVAtg1cIZN2w13CFzEN1YYCqSuQGttE1rpK3
jbxcYlee7wXgobGQ5tEPyHoQPF/74i4BFyuq98hwexJdvx9JsAj99eqCHl9yhGVredTPUC0CzGz5
bODJM4sMD+8UwezO4TsbEParofohd8VUefsMr1bJ5iXCWfQLZsB7R/y7RmFgldV0qQ4FHqbvMQj5
9uWJHkz9fP64qal+QoTgla8emfo73zUEpNzcwURruI2M6jO69YRYao28+OLbkQKi7BBBFUUe5FEl
97CGZOI63033W5JtrCvRRPfodS5BuitDs/DfK6x4GXtoF/wJ9uWxOkMtjUh51AEMH0kw/sNXASQq
7cBFC6SOUCM8KEt09wNQuJCV8opFy9qpwF+BwC2UChm3jfMW46QaNKJ7ifSTE1+SAxV3ivse3oO5
lbcte/6bs+37Vc95OAQw85XPJV6q3spsLnUK1fcqyVz43JjIXaKEj6kxFxRO7TDeBRwhQ2FiLxG5
4D6DZycBqyY1SacLkzVIPBMg5B0JQmQMxHMQSfS46erZf9tU4hexauOR3CUCZbfnRXl56lrN4l3d
WcP4Gzbe1nLfgg4mYbg38jyXpDnhQ4YeK030n5lLcSqUlf4/HXqghdCEhsyCsWefhd4yIDIhBKcR
SKdxnIzlBxJpTUAcuedCFLlb7RdwRyyz7KK7HwUBviM402wznvTCpU1q82KHYP3Vh44uX6qwU8nf
E9miL5/lyXRS/LNbU2kLZVn2S4XzD7RJTrashdClwj1jwxS03jhHOkylVdjKB/lM26rNA6MMADwV
MehIc/eGjadfHM1Ik+fYBNn//v2NtzE9XhYbakhckIeunHVHlVV9Y8c20iSruax/Nv17ygesy42G
ceepSf2rJ8BJZ17Ok5/Cyklvnx80G/Ym1s2watiIQBFbUqst58XigiuTW9HcGKgPvPOxNGvxuVBo
NVnArudt8Koi0j5Xy0K2xS+npI6J647YCeH8RfD2pfqy+Lbk8XL1cd1tl9BWxNlR0clo75KZ2qPJ
aH2TOPouSqQeoM6thvYtxcLiRE4ipFwh4vH3Ge8oUidDF89dTgaZbcHUJesEOvgCCSn5406pJBg7
AJSdKABQfCZeFsWkuQHF38sO8znn/UYtidb+P5UUeOO1q1slPS8GI0koxwWTSO4hrB0dB2erkgYA
uhRJ0OOGzsxHFWDV4LEzvz3uwsOhWepbc9P9aFPMFZAlmQ5Rq6JO4E/yEeUrhxGU/0HMeZyeJ2tC
+iU5sYkNItZtwv/BSJfCPH4t8WAWVlnWqwGytVWvLWhib9pgF2l1h60l8NrVLI12zQqhKt/370K7
FpgOElpP30XmCRl01AlOzQrjRg+ZJ6VxRbJIqEiuH0MYS9/w99lS0nlfdFH7SGA1GerF7BP5owYG
Wtav48e36FEoBH7EDxR/MdoNstYUbM1CQb1eekQNTWNEFbiwhaaYeh3aNPsw3O1We9my2gHp5ZwY
z70BbzcicvuaOF5IFafjEfq+lcWeT9D/794brr6V2N2xrcJwKHcSd8h2jdUuSC4JMAX8KCHhKpcW
rAuD8FWXlmfYJZx8VABZifo7TaqmB+ybGczE4xz4nQ/BP2742AWEOevFlsV5oXOzQ5GHSKjEtko/
p69kt4yXbR540OIAS66xkhkf2nnsYJr0XqBXJ1ZdIS4fxsBPGH3l6fKfbwT5Te1z6IpZsoC6w23D
hORRjRgoGbveoJZ5H+FeU4Dnx6SU4S+q2M9B+pCiXFQjZZ+HPshb2WxUcMC9FBs03wW4VD/u3uQd
t5i/8bjXEy53V5NKK0YNKUVdMb0SHWZY05gT2ykIFckmFz1xNNd68nvzI3oukwUzahByYQ3z1r3U
rPpf3kiFGFXhHEFyjseGbXrgCDr2nvcWM4nviltN93g2VzTuigezzLU4eVi2FNAI0oF3xu8WSjzX
qMzyl7CIVSUjn+GBukMRscGVNJU8vxcpRF1VlvzQTA5YzWPe4iMKariu/qsEtIPgUxXaECmsQ+r8
URzsRrzcOE85Dzs+G2OGflP7lLW04K4NzwQCR4Zrwe6s+k06i3vS/rr+J60iR8IYvetq3z8S4yE5
i5ZH9NtMoWbyPG1rpkOupxKwtBzut2r4lPXrI3KGWi89bpiDW/2ueS9g0QWx2CYugESQc19APjav
kOZsOdjgL6bHZ6VK5i3E9lcNBBJ/7LwYyH4zO5GUxwsg4Zfo+72rfPbYCIX6VhxfDsmZzCaj77EB
VOc/B3bnbQjCmT3vuvv9hDBzawFj+CIZv1KkCmnIRYSwEZ/17HZFldNDHY0dMcikQvHCaImJu+CR
66bu7e/ghar1hiHzVSQEo9G924p9rvhq/voWfa/7cqlPTkpMrygDv0dFR+4hnr/LAxILdT4mv0me
8fPTbjMLbmtVDxkobN7r9gNZrXzIzKfpNMdQw1Az9JijGNMDamGSDu7KoLyXmZwsiuj6HOgLhbfM
9k/za91PL6dpcUfSVM54koI54v8AfvMADDgzCp5iDcPoFWCrBAGIzB3G7Ll9WWD0WrjaQixinjMP
W06tb3Uw4y5EEJMctp6ujiY8JbekNzh8Qd+dx+DnsMb8kWHH4+2E6ap1hc1L1OZWvD0A5QybOFER
FWXd7dJ1I25VuQneBztybYjC7hvX7nfKGXlCXzU8mP0jMBZ70HjO1vLXl/HYNlFPh+ZmjGXyhLF2
TseA44gn4a333rq1Vi6cv8roHe0tAkIvbm56kKP8XDbI+yLLzRE0WKamVB4UaJ9fTBlZq30PxTkC
srzAYfkv7IBYRsdfIrz4eUEYlWQJAW8Xi5dYygd0DVGYkIrHoG+AB6J0MalBKc4E1BN/GNSeSNi8
X/pJd+L9zuYsMwedMlcnmQeDGWmEhK4+rsulNTvkx88fMTdbKT/AiYaMjF9LeuLbiil9wOGo92my
1b40kpD5EbMmwo0NJcpEooCQOR5GJbC4iVF4qePcWmyebr0Dp+uHfMNTDLS4LXCoWVhfOXAqGLjZ
ojl57crl6/jCRfw4fx0le2oiEb2JxT0Ul7Ar1OqlXXzJcE4bRg0jFjep9RWEy6drbp88LBEhSg0B
TOf77ux4kpV7udcZp7lzM+22mAdEULcI8LZau5V3MXOmxSug6jxYiZGJlJ4Q7XPvU238APCe9JHa
x2F8+IS57HU1j1UKD8qp8ZzPMIePFzgneAIcfh/pFw/V8q53kIrPkWEx7I9D0kXb0HFksRnp+065
5fvO2SC6x6MpN3DwvVrR8e6cf0+GUXdkNz5FY+u/QUgGuLVOmaMby9J5v4Wln0nDytbHJZDzdj1r
7WzzJyxSNiLDJ1l/TJtRVFp9ad/9FtuxNqzgf3krQMn+RkpFS0bVH8laSSdZYgUjB6DpGW9mMTHW
oAN67WltpHW8SpAOCeOwTvR7kAmj9gq7Xl/a2dDDZGZ5riqv1egmeEMdfziMBy/V+jWxtLgV80EZ
N+QCVH+spReGBGlG2cUpdAD3Zv9i/bleddZGd0mksbP6+yE5Q+NhikiXqr0IAdZpupMXhux7J1kg
VKnt4ainmC5VAjv5PsWPGcFrJn7aP4QSZbj2t1XGU+S6zx0V0eUXczWnt8dM0NiCRWu9zUGGlhEh
ucFnQj1mp9BIqgvvhtlq+5QIRPAKccmJO7dkZDZlbcUjAKF0s3KAZyldqdP9y2w0Y81xTnDYg+MQ
UKzBtD/zLAkbl4ViVcydT+DKmuCS0oGk5aSatTV+GnHpUnFUTss7p9M9G1wrecoltyeXPpfjpgll
zLfA8Wcwbz2SUyb7Sqxaf4ijGPJfPHj5TdEPqlj5pGyPGl/NWotIHMlTg/KBhYqhq9IIcLAbDmUm
jBsiK6pYP4nmBvLlVhXWcqTV6OyEqnx6/LPZCNxbSKayMLaaQ62yaJ0G/SwSOBI6KwiFKdYcS5/l
isvM7g87jd3yGEX3BHFCXmiFg9Wc8mwxneDPaEWjfbsHLQUtnkMQyxlPWn2l9ID1VCSkYeJfEeES
f5t2bqa3RB/0fyxaPsQXLjg8d5xFUrWAlc47t4ss4oqlIV62BJvtqtR1vJQBVde4TsqBD+ggNMY1
PGa7gouYKSs6ghJ2p34wErKiTGVoSTl1FC2n0FFv2fczlCCgpftNBS5CiaAjW6PFXGgP1rWTA+MV
M171NtLZo+fs7vFQorOT6UMeR6OphBtCfFO+W2e8th+fatJZMNyrz2FWgwuV42buxmBPP5W7YxZL
TSUpZZyX4rWqFtFXLkF+FPsw+MeHHmdD4uTVCHZNKvPPLDRw/sJP6aOGHoNCs/J75UGKTLt+rA1o
tWXBPjpWVF/r6afEfOOXt/+UnhV2Oi3l7KH52sIIyc9XEMhO0e9w9NVHU8TRGTSJoxmxAWXCNPeU
kvhb1IzTzfhRdr1Qylvr2GNapzf712R9h01JKexWhapLGS7+jgtvA/NM4z9jRE/qeJlNMafNODjo
DA6MkbgVx54lFnDvyMo1Z0lHbIFc2JiSbZGirvEMUMaEMN9gO2mktsfVdXRyc8yob36qgBAUbmiU
YvdW3YTGbF9mtTvi3Rg+wAYcpzj2b5VrOWIOHxFAADF0D0qxWtu5KfFSmfi+OUd1T1/A+ZV0jqDG
8WEffXDOvhf9pRUYltcR4GL/3JDHai66rnrJZDjCAjxwGXjYZbsGGFGLiweUyOKlXCDdemtre3y4
ENjt6WAG9A6zunZFPJuyIvz80+Iil0c4A3+vOUGOPP+zG6BIhvW3MoRUGEt1Z7QD71tPWuZKUH6T
/FPAg2+jNgfW5QMF2+pOuh+q5+gVw4ysulLJ/tvgjZcGM1ZqhxQ8rOq62F04uG80AibPY5WKyGPI
8nB3IOSkcTxo7Cl4UCVHDWvnWPhDmGmceXPRM0Je1loewK1W51TXFLjo6Q1xfSagzi+7dB7PeBds
ZOG2+IKCy5THIRJmOQMwkglo9/XsagAx6yFoVbpCifuyhUeIcibdLpdPNsIDeGYQc/TJKBCHfOuG
knhxAQp9IHRziSYTn3NFJX+AHDe+V/gwDZdPZFkccc0a+BiWWe+ggTD/c/46KQ4WZZcYElZ4B8fS
nlnvnzOG7GFa4pr6ZyzWKOiEHM5xMAhJG/95J/q3hDZeXucc1ufDC1mFJBHvvAYqp2cS46GbeT5u
ndSat594rHpAgbaQ8U62RmUoTa3UQKXoA78BMl+9IfoF9V/3az9n6l8f5vjb6FFwAfyM7FsGs0n3
5gcUFRmK0gqjG0R8CQ4q1ofrZjQgn2T4XXmYvomq2S2Ic02GZvpRCeo1/X1K9dSodalm1cQ55vEt
dDruLrH2smy+XAv9bWQ/pIuJJqwcovoxWh2d7dUc/i6Wf5BWNwM5cSuOw2t+er07R5qcJz9kH/cE
tE481oyYxdMj7ob8pRGv3OU2nXtBo+UL4cGE/bRBnvoiEArfPHRWQLUWWBl8nrm0MOPd6tIecp3U
PlFLEflM/zJpHIErL9P0SdWGZvNt/88IskRSRuDLDIzu92LILnm22i0ktbfjr7TyGqEe3WWyoYgh
6OtaObm5xYQY8yYxi2Rmxn9swXxMuN6GgychJjwNyVTGf3MV3FJkBlQxPrtUiet9O6HUZUbWlvNR
7UnkXdGDxH7Sr6bOHUtpmwcHdsTQGzJRKb7B8fISg7InNtIoiEVkcVn8q8TOrodWh6KPbF2T2WTc
UQuyMUMvjQJP5TLEqeyowymqq7HPozqkfvwe4LvkSS0a9x+YaAN0sUhbwf+xCNZMv2hr1M6kzvD3
2bAzGaOX7PoVcOdGjpJ86g4G0YJ6vhRzZ/oO1+t0P3y+i+wIIJVd+HwFg9kH4n8iYvophhf9h2rE
8KZx8w07nOEbc/7tbwCA/770DbyA0tspZiD3OMRWuUgyiIBkmhIP+2m+VeeLqaVoW8fsdQO6WxBh
oD0/cHlIep0v503+fVvEdDiVxLQy9i+zxG02N+J3qp/2nXjOrC+8TdYy0cw7tqnKnnIZSgI1fYSH
3tTLatS9b8UwDK6SmwPlnppDu1E7E3YA1oTi/kZhsdetCZNa3gtygtvKWWzx9hu1oq/Aa5CbAe/1
TU8QyS5zwOk3omnuKBla6I3GdwHlfSxAECLnoCOrpebICrcApuYyBH/Ehq/STEli+LhVSUBrEacg
PyzQzgDeXYwH8ei/udq4to9eSXdBy7I5+xkXUdf6HtgHysAh4hQl2LNgYvLk4zEsIGJr3a9FNFkF
oXjZgc+aIrLJkL+a5ZtXSKwGluugry+Y5XDVnTMDhWmZmlUhsv94JjZq3NER7rKSWQiSVAOAwb5W
FTXgPcJ65vp0ZOgCJzk1FisZBoQoB3neRzp+fV5USyGIec60KdgcAHT0reDtns1GFuTJpRzfUnpm
lRWk+nBLT4OkCtoWxgKf2q0JAn3VrFEdqI64ARZB1dM2aARgeML3FzKQItbmZBqUtcduDCqn9DlS
/eJ78jXp+i9+wUvSFuWcOecyEkLkCmyFzvyTP/TlouAK13n6aQpokMaXfWC/ewLrlisITNfg6N1e
9N5IbzRf3a3k0eotLAsi+EOJQeZc6u1TguRD/url7aJF2wL/hfGx6+dt7/Zb/T7D/2DAhfhw0VQD
ujUS89klZSstcrhmacSxGJNof/ksPjjr5dGi5g6gXCkCMVLoHVoSyIy8oMF6WPSYD6TMdG16q1qT
fsoUylm4wPiq958/ULiGUf8easv5QC/8Qst4i7DVXbOEdP+CczG/p0mhYTLf8/y9rRCvx6s3tqiy
IiN+0ldEXhcg+C0V4wjd00EqFu9+Pdx469qHsI4bi3Xm+pwdRzLm9ec3OYLIklEKZjnRfkbWT6O8
B7Llgs+dR4821CqnZF57z1ndOi0BiOYMKqogoN7tZaIaDufICTlmUf8ldYKBiulYm0Yg14Nnzakf
H9Wp6rscIplzmPBpV18Cl9UshTIENLRaMHU4FWWeBzAWUFKIWcxrPNJOpM1UvKvL+PuqjsPLcdzv
PHhPjD3X1FZ835tn/eLXoPr3OlertVIU/GLg5dWdNpLaMvfORzZcgZCbVnha7CTD+3zA/gW+opD9
IrySogJScZ3Q+rsE0W7f5z32JcdDc9KkkNfdJt2TRUlP+Ok034m8JXL7U5jLx59Vr4I6NjOhy8O5
h5CxHKrPsshrCRqeTE6vjduiWdem7y+5GB8dbPs4bBr4GLc6yr+AKwASqQNb0ZdUUSZEM7/NSgbQ
S6jojJcPyPdPtnjFHHEi71msylPzCnpGSXhQY0Wf2sV+STymOX/QtBeDv8McmEHdytZKnG8l9zxB
baxdDCpL98FOLB+h8W1LQd+2ev9a01ijtMNulps/EuVk0bX7KzuR8aHyZQFcsN78Dvpt9uti5bdR
0EWOh85EvZlGv/Tz4xBdzfhgoX/jKKSpfxMO3DG6p6c/QSBALmNKQtXh7veKqZZHlkmvOKMBCLUD
D4nKhT97AZHdWNYhI98CFNmtNbVzfcxoAWSVa9n8VSTsxa96O6IWsscICg2FjF6PDFBMFgAfqMUU
2+89ioSUiej8jdvCOcOSuTONYSuz7ShuljL/IBPJgLiQ8cOo030faKK3EAhyLgp3Ydpod0klMpRQ
5XCggbR8OQo5jATNT3S0iEwaOZn19Jyy723XpKgLtRQzAWV6lBf4dojMl8WfNpLRDMWOaTSAHGmI
JEaXYVaZSPpXjwOMQCaXhIWLqkgD7LxAYUA0w1O7a1sE2F4xuxnK3cEboK79PRT8FO0XDzCjrhnn
irZ5Rp4nWNxqbBV3J5le3Kv+h7ASmz2ptHN9rtR5lUNs7D7NvgN/ARSYTAqrOUk+K2KF/1zH+u9O
uVPDQYvn4k+TBJHM0M6RD7+R3hwMv3i+2HrnTnDxtoGbO+8pU53MtZlxoKYiiGNNLDmXHFFlO8Ap
5DbRoqJrarD62iXigSOyqdQ+jI5QfZzEuyxJozh3g1oKDFFP21xURsw4QaVOXbZVc9McyHifZp4d
e+IsFLxMmUTKrNhGmeFBpN/VFIrGuBGdRZJFaEGjI31SJLDzAXPin0/ABaK6C9HsKrD+SNoP1OoQ
AFlvZikzSJOca3Xj3/Bn8rBvW24kdve1Xqh4pFoC0uVbO4AHJkirawJdBJJVGwwHgmhlnvaU2nQd
HqSlpZEUvE+c5JY2GKEpLixe916XzHnbJR2VmQxKx4XTwbedDd9Rdsrg/Znuf2AjWPhc5H7JRdok
k24oEJ/v2AvrSW4hr9MK5LsAXCI5m6Vunk0dIwP+ueQomM+Bstcf/zH35VJShI1vE2r7DIX/E/gd
teJ5LYKxJ5ZOcxIJWMxHUPwB9x4T/sX7QodEKjSPAXPx5VoVT6LfOAwGA8p8lsTfHbCl6wKkokkr
HnaLfpCH42vGj2BBvV4St08is6roR+SlR5/6+/LwdJMZoy0wCpSwej0ni82YERfB2I8UNZxwiDV4
LsVHA4FoFOgKAV7d9L1rpn/Ug8zurnPpLHkxFYO/gc6wA2RWuukP4tPyjdp1MtZ9ZO/JrDyrq8ge
BmHaTY4d2ireTX5BvBajARvSfm5Y+lqou9pqblkS69wdDOCFRiQ5Tcnne5wUC/56qxQ4RJMrnStH
9dtlfxgGeMjuwE/RcVU4ClWVvsYd19j0OjDM6fZjffQxWxpgtkjzOF58HkGt8OfgC4tYmb2+p7KG
GtAXT0tG9Rcnt02OViOd3hlGVXOxotAMHhJn2KqV4ckq6ByMfUsAa1xLeFkD98889AKMVnx4I6B0
7mBS6U0/8GfUi3VSlxn1uv3qK+cEaxlo1gkRDQGQTrzL6OjdhLxoOoOxG63PpCqchPHHNJaIUl/S
wP4ucS+t+0oBb/Gkl/CivL4eEgnehqxz8xQttVspcTNb/9LR4fpcDA3GIrDoQen+DjHdkNJ53ssE
H7jfOC/4nCzf0XwlAprC0LAvxDH/B7rzy8UKE0GmTuMAzg110s4ntObmjav71ze4p9Jmn9Z4KkeK
3BvDrV2A41pw28TD7ZL73Ht89X4NcLnjjDtgMdQs5WtqMptf5kpnNrLsWJu4lzJWRKnpuxctNDVp
KaL0niz7Yj/4UskrUksUqe2WXcTX2C4XbB/oZWvfbUu2HrC8O6f7otxdlcWibgzWaLnpWGRsoZw0
wCY+z6a5WrQ8yTzBMFDCu2OPs48asjig5Zr7usoyzWrMjAVZsq9BtIHzuVHJNFG5i99suNLDORXp
10wZV74ZYuIf/rLdbxc4m8u+pGMyufi4IDCZCHXK1QYIvklvtH0QkRMmSRej85B+2DmncxBCXDPJ
UBGCdyhmL3bJKzHhdlPirSZ7rJKwhwW+AxTwRgw1OemIMrZjeZNb7xB89YHu9niQRbsv3uE4dMMG
YGVYOKyRwAI4M4rOpHgsnuVC5B9Bl3QsWHyZnEmp1qKFmn9IHjVDaxAB4xnAs9esLFRQ9WgpFX0E
hoNG4WmOyYlfdMxnjKQvps7IBAUn0YcxGcPfeyOCUV4aihdFTmivMJ78EuvMe7xZnd4JmHU+CJ9J
yoUFoJG/AMKqa13fQwSY3OvAaDWTZ5Nw0BhXQ9zrksGve781314XkiArccYyr9D7QHwG4LNGD8QU
18btr+Cr+ikcxs/EDUQSXfUpzYAygMHN4Dk/DQADxxl6y2Hmon/NzeguAv64B+9d3lstYmTopvMc
E7W/ljYrCjaNu441i4Qv9e8wkbmuWLIPR2shKD+vaMbI2S9jVBW8iwqGsCcO7RdxRrHCuLceCIUf
OFXXqA5oSscTnKsvpXu0R5U+4BVY2sKfsOwEQf/gDzZYGoQaIDMRUVxQD/eDJQnUva4VXQUNmfEo
T+gpKHc6Y3JfCgXQ0tkN/O7TUbNQcDDnynLf07gvqe1dY6Bgj0L2+awhZZasqmfHse3YntPoWW7O
VvqPEV+ClNfzVNFqyhPrIuowzBvb//D64+QrS+eko+zF9RI1mQydLwLcIP06V7qGAqPNl/H+ZK4m
eXpELFrhvTSzYDi1p0NJ4DUHkmNA3z6BmoVTdYV+vHtPWE2JfO+gd5NX+oBw5SS912AanIARdPVb
QV9YtCzKDaQapQEU565LLnO9XfXgWSObdbS18+4zfMgLLW5H7FN35p26Xn++hTEEL0qFBqTHoNCC
dWlT4pLeulb00dKhnRQAXGa0tMRWfyc5XM7dCQDOWSRFibINVdyrSz/5hb23t0RKEz3GvOy8rzPi
NXmDXllErtd5EkS1TA0adD+v1C6vOAqnqoZH17wocwOyB821v/OQ+qO4NwzMAXQJvNU4W2mn0SGf
lbzQg5m5XfCXjAC4brf7tAPi1C/MZx//r1fhCW++L6zi2dYBrCx922T8AfsfVyD8xfkp9PyPkHCv
+cwWvfoPIjCGJGsJrj6HOiIUnCXoIDNaNbRipMK3fqb6MJtSsj2N/tblnwG5JbVgag6a80yYk5Sd
I723L/vhPafkH93BmH33YHJ9knnd9NIj6Jgt/AafugoqzJnvT27hnrNfjV4N9CB1cBFn+4yVrQHz
HExx1MmitiK8BDj2EXs/Jp0E3bMOw6oCy05SwP/EFHfpGHKNSLVhnQD71IS9yyXBDYp6B7RNS/3b
PIAKRuCm7DJpmdyCmxvQv3FVT4gI37wr29GO5BY3XL7c5foSyUIlKMgAPPxzvgmVC7L3CUaBkE+z
omCau00kvpm9B2nRB/IszWPRYMycBMxlRtIAgXoqEyICd2qF/7sh8fkQ3+l3C9IBh9HFBmHEy5h/
cRDbYP6S0TJJQtfpAGAhg1KqWUPdm0qdSY8mHASzSwzfr2yIyni1rwbAXdYSHr8OCj/RwOX0T7kc
CZek+DcKEzfSiwAu/n+UaoluE7ehXmwLm8t0V61fA9a7e3cnerw1uDnn3OKsbXQ104RI41O+zOza
VATGTDQHTYVjfrVt4pWnqBdP/MDPYop07XIg9JgWGLCXOlLcvM46VMceAiAvLB1hH+gkoyZAqA5M
uVNnT+9LnBtuybhKR4QK57+XEX1POpFuJpRx3BUzF+XlCoFNMXprk8JCyjDpTr1sE7+Qi+J9IGGM
2jo4UoERrOFaAgUL2s6CYOnADJUf26AcYtynpckzmlz/rD4l43/VXelEpGrcM18Y41TvodoLB8jN
G8waDhu1VX+v5JvHiGdAVPjZ8wskYWO6U6HFYNEwTfhTtx+Wmnp4jmvyucMoyc3FOUer0kswrMxC
2P16pJ680qVMYVJ5/VUxTJ7UYroaVxeIUF7SuSpa3dZQlfU50RuUsotemRaB4r9mu/dvPQsgloNx
wUa4dcmZldwHHtVGmDCQfRnu2CRkE10m8VHr9CQqGUMykeUromdQNYEWXQ6kX3pvw7t6OXV/cuce
chJUV6c4SGl2TKxUykSuvLeNC7CYd1idAxH9pBUdyOu5UoMTpuiaChEM8j51ZveJrOqdnQsRnO1D
C3EWWUjXx+SMCzodhmbyq+eXo1HjRSpiATA2nGr2W//R8VSbTz51Tiugz6uyu+kkudxjgsJ+iQRN
16x4g5DbtpmFO3kDVXpmDNBkp9QVWL4MTu7V+mj54gg89Y3MBsnigfzGe1tlUWK1U6M5TJrwHbp1
lYYcF6d9/aVAfrqYaZM2NJs8Pftn0q5GWn5LX2+cd4ZRGY9MN5oNL8L1Ctnd316VtqVAhCP3y1v2
elOioHzAy1HWoMllnPhs7bpb01/NMS2CgiRXr+IUWRdas/t49WLhtftxoX6qyepLSjZ3a7zw1dbE
PVX3+w2g3DqeuRE2Zuv4kun6SrQ87dFmN4bf2XljOf0lfx1qT6ceOw8SkBtQ0QjoLmbtwujpBN3L
d0KJMGsoRNqrAadSij8i/35MK0QnCCTgxTVN1hB443Irm5qERpoyV5fh27ay8Hocemvr6BSThzQY
3RlOsYlubiy4w3/QUyjVOBy4iVJh1cd4yXqf0YkBRKlMP4hN++0osV8Y5qP/QHGBP0NSzkBeRZ8K
Psci4evGjJuwr8Vjxig2d3yKfEmi3KK4ixGM6PKrrapLkDNzITEO+4OtyQnW0j+M2lL+KZglzwZ0
are+QSnrnTZ2rWEvTLfhn8quOLZMJcEpSRznSysybJ0f8p+jI8uAp7zIy0b0PA8eFMvd0BFFiqN4
ooDJRJS2f5X6KOY2jWVxQHQwssZIIdcQLzIPNkwxVUOuxrrR1DXAY9+JvQS0LmsBtsRmMn65ET5M
VZga2ZdGArmbpwI6s0+dol464P9pvnrzuxWzwLMfWOfs6gpOEdrfy5ckpQkcE0KEWi7+Ev3BFUf/
ooKTtX7LsPzIXl4xSUzH69+LDv8/jvvyc08SukS+vwygChUhAtYZNrYMJJse3RibcQjEQokgshru
V9gx2AQ8wKvtfcUPkFsOlQt57NgIGF8AZnExFpawSz7iKEIZ7LQHtHriqnrH2UkxQ+k+q3fL80p+
kkIzaWz3FoJj+GxvHLx/FQEMAim4XKCR31UhAzcPQhzbynbXqlWBgcwPJ/fWto467Dc4ZTwrK3GO
aFA+4pTKOhqFwc8T5am3VMCaWO+gDXaU7A9zbLtZK1eYo1mplY6FcQFnUs/NMdR1Hj0r5WktC6uB
mHC4leQdL+yfsrm4zXQTP7h2zVmMZGwlFTQgPcuXYoxa2IKm/YAsN00EL9byptuX9H4P1tHl04Qn
AZ+egsSTGalyhWnNgtWqM9UhqdlzhZxNMalkWHvY/CZnjWUridRWLeptBsfpj/zoaQE4FuD9vCBP
RyuTOhHOPq33PJBSpVVLOt0gQgVBgxPt35YLC7zdowBGyNEtt2UZTjnZcPKWpq8gpoLxSyBaoKFq
55PquDXdkq+ztOefz9l4jmk6IqPFuTz7UW5DI6Org3/M5RG47E5AK/C7jvGuWIXtGDRe8QzE/9WF
J4fFzRvWpGyoAp4gn94VkJAbxw1797n7AZOF1NAFM0qj4JXtztokdhgwHXUXl/JLYfyjKQBtrqr1
SHQiJuhA/VEEz1iT/RmstNbvGOsTdRCFWFjTMAXU7RUtCTZTeXHNS2LCEZecRvgWl63MmKEPVvox
UiA5KroUxye5CbuTIFefHByRHsFjbC5Kxu2GbgM9VgF4BNJaJGJn3w0ITAH3XkGIqrjxlz05NJyx
6BqhIFSJ1ozlQFQ3XKnd0X3pw2M781N357qaxIQLeTvmLAAGHqvMgjXKm8umGK2YJ/uvVUyVdRXt
jo0rGujvNpEXEYOb2NBp4f+7DXYsiafVqOivkdAi9oulqjAqlDalwzd9qXrbC4PaYNzdzM0Cn0xP
7NuQD0C3KEZQc1lzjyvwiJa8VSsUPbThKUILG39RZC67daXL4svJIlo4AyxUrsYNvng5FbKl5r+C
/yjwG7GweCTcUxe2vzkgr8ijVC7cVNu0GS3tVgGZALen5sOwJuqfYAoDEsLLFRyR5NTeZxQZw4ub
6iSmkLy9oNWLBmHwZQlefj2ElJuK/H8p7HEjcPD+rWf/pBANFVLVCie2ccyJ0nhiKuYx+CTmgbGk
4b2CZaa+PEzA6Gmg+vjGNqCZI7rMuQ7mGzaRSVXS+Nxj94RVzAn4PDTzI51F72jJimcxGAYVdIlx
LFxeR27Iw8da2F4Xqi/JGPs3j4j4M0k43coQbRVZfioAaMLfLk3i8QyXrmgwACEyoBqrm1D24VLx
4Gr05/GVUx7b+zjKYGESkV4vMYvjVtl9bLcdx6t02UmBMa2j+eeWg0z/FPkRGSGptJadw3xSC7lR
fUzjCfKEla1R8vaUWzajv2scKMwulkOSdMlgx3Sr1seLqJQUqNZFHNMfOOOkFq6hXafEQ8gT+FLy
7slWc1yzjXPouyYWijiMvou+JoxKUZmWsMwe05qlZ1QAN6WJcHSAdUy0PTBxV6SwXGzXEhFMd6hB
43MMxIpxV5YRl6OwbrDypkJ2S2Dj5qA8vFjBUmlpBfFeluUJ38jh/ereW7vpxesCLqR07xXTGoxh
xuvSWKhg1Pf0CIh24EYdGYRNHDehAat2cp2fZpvjGZreIYeb4OuSFWE6/7h12H3j6hbIbJSXC2f7
ouN7sxDpJU5+693Vzt8tMxtus1Duvyo2kHNg9XhzCTA7PMIDfbb0yMnl8bJC/YmZUwGAADYsebbY
c17SPkAAvI9wsWlZUsjkCx6v5jWdIKJywmpeK1qKwAEZxPinDqGdrl9qmb1PM6Wi4o5hufjiHbwM
Ur3lLrniaoYL6Q+xll+b+zRHdckcQ/QLmKwJjm8JCznw+AI947MyJFx+DTvykQZZFHZ9KLsfKFXU
+0nsvBHu6k171tsYJlIPFqoG7AaWZK0ITqRLKuXVN8NUsBMS9ZmAt1DhMcSOVurSFpmvXVe4PGy7
CIWy0Zn7G0RVt68kILOR33/2DLP5xU6JkgXSIiWuqGSr3K/3JQmfyEqW0GVExnGej4qpx+AW1y5W
ELuih9pKQquzq8cmTI/prTgVDKBD7ZpbJJW5Ji+IAovADLqqVxnwsbBuDbGLC1fdVXaDix1UP0/l
Fj+bTrYbfAt7T2bYTIsM5zWdS0JkbcZdS4LEiFTE62y/HJLBKDR8GtrbQ6FWApFZtElDM+3Bd1Nl
lYvSWV/npAJWBoE0dFUz0ZuI7GNqeY2O04j1cgUNLa1gMWo+1rYjWMrZfeFGRSNCXTelsj3A+Hdt
qYaYapye0sG/W8lgSK127L9tGQQlH3iC0FrLlS/XkrBZ7iTGAHxU7X4FbrBsnTJp2//S4ngrM8f0
CqRxz9b6+HHtYeeObrn1w3PLQ6FQ3kRozkSuU6DwpIfOlR3NSUHyWwSEJNYQkZyVU7Je+oNDY/Md
G0R0eItJXd8ue+iMCKCR38F21wiMZKWNmRYytY8cvPu4FNORzSNwO9cNO3ekKpRTPiKbhJh8KnfW
lr0kkW+Md6fmaxK7Jtwr/nTRrrtWO/Z75wHeaxdTxIeBCVom7F/y8ad8+bD99/NEazXVmxqHD28N
WXSpYafyW0yYUyj8V9x2TpZnp9F7aH9/i7EqIcyx4OLDOs1om7KeHAQsLHD4N7AaMNnCrw4bt5ho
4K65i7Q+QkXXI7cv8KEoRKjvF7qxNibXk/BRQM5M/Vuy2pFRE7osEAq4Zuo+K85Y6s4U9pQm3xGW
1C2F/HhI1pzoou0zO/Q9L+SSnbzQRShXwdyvPvimN1DU3BDsR6bT90TuhSjru81hs/FvKjyhvt1w
D+ZRa+0b0WueAkyuRxul8xaaW54ykvs1Vlwxu43vrGJrBO08zGOvasYSzSqW0hF1hFb62/8Yzn+S
89yMCiwFRdy6BAG/GSTbKX7E8sx0azdW0PyAPP4xoYzwHAL84b8nn1AANGPgvVbzCxTXIm5pvLk1
Un8cKdo6gQgW8jFkn/1duCdkg5Lea1rX2IUJz6tf8qWytVax8Exkk9AL8zBZtipgJA3raMjnaTu7
CebelD/M5xIieKglTNrvMNP9GxhKx2LTfHSEQOXrC39Q/1rJ4sztU+yDXJEBEWyxo0V+arpQ/P7B
gIZr31dhiGfxSHcGULVe2cYRb8iYdNXc89xDtzl86XXcv/EJnihBb4Cqtc4YsCYBUD1TZR15KaZ2
5pmLl3TkPFvLEtC0dpMSt4qxMW0DKB3HZyTO45MovcJ2Y1ap8tt7FqPbbrSyOMpdQoXY/cBK7sWz
FtDj1Cz5cpsg4j7/j4NfGT3FIqQMag0zPjS0YW0BIxL+eDEOlvr9IL0NXBZJ8/4bq5OlTc6ZkBYZ
g/n5BsmNXE7AzSjSQAKRL/nLMcH/993BNz5LOvdtbzd75rOUs5WQ/DPL29Bc/mpWs4tqv92w8b9B
x5bJb+ctpmvpdSLb7xQ5P5A6x9JGDTP4C27k9VXiId/iyC7iMeCakiwTiiop3Sk4A7oqXKDnjeXV
e4eTKYrA4hc3sP3oN1sf6e8XB7zAla7rZigHPEF1lJGHhuw0EYzkp54bprHuNEIK3qghuggU7sN/
KeLkaVXhLx5ewhaUezT3sOmG+K3xnIO25wygUoUhj4HSk9BZBqJr9XrhFvzEgQCAAKTr+7KyC1nj
SigFZhYjO0jaTXMjidR9ON5NQXeIg2fmhhMgYeZeb9vaDptKdKS4fctp/hEFzlhfgWAZsKrpjH6H
/ZELsHqZcNAdXiGC2+9mDTaQ5tVOXU0jbkYV76XcwRS2tSX7NvOECDekGvPTYBPXgrlr+LmPvq2s
p6DK1175JAcLwiEVf0/KKgcf69NAEQHoTtBkHXv5f8cm+GhmUOczA01A2iUAJI0h3yivF735L1a5
U6m8gTzLKIH/CdrQ64Gd0Ddw0fapRRtd3O9abkSS3xFtDCvSbiYnN2F40XU70sFzLwE79RpArSP8
0Qu/+FX8dnX227JyGB1tnZTBkgcfk5S/kC+OgA3lChTeQ7PLlwM3LjlVn55hTT6tsZLtr8yiJv4U
RgeHJ8enOLn1Hal2ip4R/yQSbseZ4H+JQGfQaA8c0zl+B+VWZ7kl5Sl4zcCVflF6STyTIRdOBLYY
2K7dccOWQtZN3ubGFyLGDoIuKUUGzQNcD8B15eMTuJsDVexT65HmrKkql0O+WBfTl6H+0acQFSTE
tVbLROC+M6QpKzBzZ0pfeIfnmxbmZeIHt2efs/3tz4FyjCjR8rrWBRI6Zk1AC3ceLEpX4JZTjH3w
7dNb0dTdRzAWiLNvfWGrVlC1eun9xJF5TzImCCzQy+2kJQwvGg0qRs+2c4OtcqMZ38YnU3Rb+LpK
rEJqWmblD6sg2jNY0aZu+WK7amFPM0cbixOwBL55Z5Hy91eQsNYHGopfI8oZBkBX8J1wMWxmW2Jw
iSSNM3pb2OJVJPzF40kDi/OIndb0c0amCkkIjpcxggjPlp9has5FZ+g5cKmaR28kVGoDnbMsVeO4
waTDksom9YXW8S01du1laBFcr6YBdqLc45qpAl63JHbC9Kew0HqeHXLKueIPh2JodxYHTAnt+QBV
g189yeGEwiN1Tf+XMzDXSFZhf3ZJljtX9DpJT+EzoSj1n14aisKApZ4nVX1z8YjMM6wPmK9KBg6/
8nBJKGLIbbDlPQ5iCoKH2Wgv2gwdbWeyK5KmE18v7XroIf0WuOAEYRlmBa61Mswd5T2x+kfmGyW8
1BrZxdl2kOoV2xMXLcQQUETTCxOqy+fSZd/QclJ3pZ/PYCpoYKdmOda7fMIrCX659f1FM5o4VTN2
8QzW3CG+QNWqy2yJfILtRwJE5Wrak9Uzaa2iakFd2gLCpAUlHcBlRBDswtmeiB5sy+4KD4zkNkac
CMoIj3qbhAqxwO0Ks/Xr1hCEUpIJoE58sg/5o7LiM/+S9Ma1LqybVbfxUt5kf27qBTj4IGwSGFJ9
puMrghtxd6y9lCwQajqCPU6NT0Nm//PCT7qO2Bhy76OgT+CcEij5XMU5FezTs0nhSPjc0Fcbsg6m
39uGz5XVUzlwdDVMZKnZ5i++iSojGn/Fa+V2MwqboTrkJdPxum6iBOkW4Ey/4d4O96Wdm2QkCVaX
3oBRLXXodemwTw9JYO/Qm0nhOhRvsQic6LBVVTK5amU6NF5j4Q5XyqwflSmR8XxuSEXtYqDjMmzX
II/RrhImpPfV8nXlr4ka6uXi2ZmsF/dcOUa9MAPyAkIvFi04DW0x13gWHx5rXDT/u2YExUEOmZBg
T7cxI/pNvopYjwV5yrFQIORUiDfWTg0e0eEltmM9FOBlDBwcCVfDyQVj2zDNH7mXAOr8FnH3dm6n
UbpiDVlOyZpzvPr7Up4W1H7tHNNRmftriSpgxf2R4A5L5ELtEfUtHbSylqiRJAEIE2/SMipV0zgV
NluZ5c8jqem5DYZ55HWzYGxehH5RhUJPqSyj00uJ/uK2HQWJ0xRZnWTZyhMmHlsTxXFZ+8mtvZmI
/V+908RcqObjAwu4J+ypogaM5Kii3JYTJdVl5RtLlrCLKy1faopZiVbBxGfAUO6mazawAWi7dWcc
0/PfLHM/3+mp8bhA86JX6biXDIiXGVlxTFeds4ErqSBTU9xqZDjguHa9bgoYY5RZul7fibDVLjtF
DyHHmo2/bYfuEeSmADnTZmLYcVVlhRAhikQQSZMQwWRmkw6qEnXgDRv9cCtZt0S/KlVPEoB6jj4h
PeXKD7KYDCHM9soZWoQNE9uSa66517LpYfwrC19hhpl8XkY8w0Wu3RqSU/mpNGYoWBs0OO/UhXQf
BgngSzL7FDuOSSrtpNbbY6tTZZJS3QQez7RSLY6EDXxxvhEe+bNEJg6KS4PdsfQzOa0xbTQPxqiw
rk+5yFvEWiwwBPUcbq/XayJ4UiDCzYlGTebfIgE1Cf3TerJ+oAf0PTSUx9si99uIvt16S4zYIgEE
urvpBgcBRUo9nzknly4Qp7lkwE+cAkjLCPpqpLAGNot3saOsrQ+rlQk/W4tIx0s37gGWi2uWDN3u
WJgs9RXjqd56ejzfcMwuFjWRymh0ve9hYcaEsO1qm5Dy7N9wwo9s32m+4FeK/e0oTrVLk1Lb73y3
sDdldW5Bl+5J4kK5ttGrhWOYUOnIuIASAMkR/NZZqxyFvQhEgmx07x8M8fr/tPuvLdx1HOocPM5s
K9LGbB9sOzaDyrsvqZmOo9ki2Y+P/Y6PCk7mjXs0nAGPe6EwD/c8ghRf8wDo4Pn6T+KAtQPMQOdD
+rysEjgxHgPWAtPj0PDtbQWAIOaSR6fLycag+kNdZm/tllwmMDHRKUo5ZZHXBAkZd2y5077dcY9N
f6cGZgFbgU+8pVzT2d4HzIPIhw3vK2JrWy7t9Bxip2F8gqJJ2wA0rRoviwUUsVBY9rBofsHfk32U
dAvq3BRZb+PvjnrFb/Crs+WrE15QHBgSoMKIkMCxPLkdpj5cZFhxeGZwAtRgFSwSSIx5e3Htbmrb
S6dSeiaFtcUTUomK45hkk7qPNdoh9D4y3V8rwpRlReylX5Ij3VvJLoEQeDPe6n9UWooBMhJG4/dC
A03JdgD1f0VLQM3vCtMscociGQrh4rbU8z9oBUhLGYZx9F8VfsOEm8Gr+as7JyQq2FDwe1Ni+Nhc
Lgbx5VvUR59+jPuEXkb6cNDPeclvOj0YMYhu0/Eu5hs4OZjezarPYtLKeQp/i6mplU0sTkEew3Xi
kXgB27/u97daFZ4j20rquZLZPfNemSbWQLMiZxpiyPQRk64iNTzjrLqeeR0z6OwusUJ7dOzntGJ+
vx3orhg5Rmz1NTELK5FU++P9eQx2hzL5s1uzwVyS2ecSHPHkO1ruVbJGse3iy6oV0uS0wpU+mCgC
btqIx12wOtUnlFRGQqljGiLZV/pmHowtJKV1RpaJOv6mFIVXtC/Smzh1oWeaEbsla45nQuq0AwaP
+eBc/tjn2IsbrFO+/mR3a7vOHwYlFOStwDjqiN/E+mNKW/cb2Q93wdDwocnLwCxgIpOmVTDzqELl
xSR47FHEb6VdI9YXm3QysGEpU1MMZ+11LWlAXLx5rQbj83l4h/gziHfXuC++xZFpNWsYgngJOYE7
d+Nbj8HqktvgnZ3cq+zIgqLCNdTJlG9X0IuXgo6whtAgAibaHlDjc5xHq4nQEq2InpjIzBkTfczc
y/NjLxnPR2RNVquSOPo3JOUOdja6X0cIGeV3jk0BjS2FTOsa0oWalea6Twbe/D2e/HXv2W3wuQuE
ouSbs8es0irZrLDwVERR3ftp0N46iAbavbXy+qXSYBO3HPLpSuZ4P76tguut/4BdV/kIPOXWvgbf
owxctfp0hN8UCkzYECOkakVfCDCRjVHGV8bHvZyqf+1auylkcwde9mzgNNYIDz2e2fHEIgbeK7us
u+u1zcdZ2cE965YIeqEUinNigJpcpBUcQ1wC7lxwfRgp/vu6owLUkOZpQEIa9jl/0Iw88ZD0nfmw
xyXRc5igRrlfeV6UKNSal4x+ngAEz+DLJdNK10YzM+vZRWrlGfQAzhGGuvT1mn5bpN3ez7OmJqJd
yjCxwaGYPxZJs57sHC1/wi+F293T0rfcstY4enrif8TrOdrui8lIyS4q9Njg+7boF/idU40eB3an
2medVURr2hPDFBztINLyyP+TZGNt9uro637gdC4BmQWWhGBeciOUXDclkkIs529egtMnv3yWKrzQ
Icv5C37ad0QhvP1N6S1R9W3OB1qk3pEUwtwDUCsQe/EJrntbaIgNoRPoEx5Hti81sWv41WJx3W8i
kbVzazlB+Crif4tmdCczlTGBk2FTq+24axI7iqMV/33o8h+TCTjfvYScHPUq0kH4G3ecbYCZrd8j
NltyaRgmPxmc6l41Dhy2Uufw69lo3me/tc+B61gbc9FLtLh8G9o05J8/LO5YD43GNWMrKw6Tiyeu
UUnqVueRn9uyWNLjtLxXnjkNB7V5ihpQUZtVLZMI728z/6eityR1Iufv7fXrTOSUv5lIru3C8c14
BBLVwo+952iIpKgLWdq3VBbmJae0HWLV1nrVmnQv7X3nBHTvPDbzBNkrhWj3UBfq4aH+NtMgGTOI
oJ4WjRMpoNkthMEy3vkFwwn54xTNyiuVi7u25a22gOSU/QD2TcGI9/sb4xEypixoTGM5Ps0nqe7O
JQOgE2z1lhl1lI+z0QAwcJ5j0aoNLm8m3VjbtvnoyrDZbW6tcpdcFvvno1YLJU5shNepZWxAcHuk
ifbeTeRZ5+LZXcR37b8CIsGWdITpbwsC5EbE7T1V3UaQN7AoL05BD6zKo0PVaqcXUq+66Z233Scz
1yNfeLwQPb/nTOOArwJSXrRUoR0KQRIklSmSbp3nfC+JcNBwNxLzwk2JOGC0QOVMDXGIhFZaKNOd
AykWgo8FFrSaNqnV68nN7Wh2UqDWP5RsaKyrMAMqrgtkXWmys7mUkMBAayNG2IbkrMXb6NFWETG4
fEZlI1mDFv+r+sc8FgBEqPjIwaDRKYyuhyT3lXzKEikGRpuXmUrJgAjE80PuupxQlGF9EbOopptN
1M62Y4GPo92oQ9bMcJFExiZ8qsj3ZNsJTgJdKp0Suwy3t3iF6vxPJvbU3ZhshXxjyHnAsgVo637f
yKdDiaz+UShpR2XjW4RpauC4cAdFTtH53B9qmWgoYKLOiBmGPxGHieOwtN5wr7pxYtTCUmqVZxgu
HKd56aB3dAx7gLb7wj47x1c6mEJVg2ntCano1r2vjMqwZ02VCp77ixOpYr+JIxgT+EpIwNykwYxC
kVZTU+m7C7waMV9aN8CsAWLgCF3g8bYJfVO3dDpVRhPH2VsKT2Il6vDlVexN75Ns1juj20EU85EC
XCCv1B94oEewAtDKD8cqfJ8I0yPjYCMR2gIZ4UGOZIK5X5JdgedvRlZP8f8g9JGjJbxafyPKf6Mk
cHVSSQeXuBTUy+dYAtfr1edIpyOwl7ptcheoA1eT5OuWnef5ZRUsmGqG8KivCCtmSA1VIoP4XG6J
+KwjS4Z9QG3PTOn7aMtZou/pTOBGE0PORGR657IEN3MPo/YNO7yoStrbLZn/KmJ+cT2DDDy0OuC+
F9QGWiLY2LYNj0MCZDP1gCyWRCetgE2hGUG9CY2bOgA3c1e4g1PIA1yjBt2n+3Ulrr3dAztBZdVc
xE3X+Ktyj/FRr6cKb0dInhI0ymNxhkvyQveduK/gvGXHDWBtLLH57CLav3uIsPLsm3ICXIkIKnYh
7dBjxPksFNzeh0gYw8bcOqMvtKteuyK822VHDDL20oge1kI3uEOC/fqorFWinzchNvIi+zfmhYd5
yO9vbxS/7KWBFqAnzllHWX40znpruLBORTBpOQKHbQA1vV4qmSbiWqjOwW0FWrZ6z2N3Hz+Ibgo7
Q34+yN7UdEst/aY9jh1GKIOEA5a35LW2ilQW+vEPWLTMwtSButlEIAAjbAcSWme0q6xxJKDenk8e
+gWys+Gb3vijVTlCQzQDGQGAuzMVcn/VBBcG4cmVgrMJxUVBoTYBSu1YhL62ILD2ibvx/+Jl4Nkc
tgzFpEEdzxalCeRyL63+2NwZnllHO+HmRDGFibwkVNuxeuSl5q3dvGNf+uTCBDUWR3NWDZ+m/mK6
MwDbgEcWvX+oQ3EuTGXgaOUgZ/4LMHe1RNNJk4i51jTfQQsJpUIwt0KcOqZ8t30juUnVytizfprr
w4xQLPopQQZHohZAoBK0UNPTp0BdiiEI57mZrf+0miFxzCIaCPubazp922A+TXOW7T008RV7CwLz
WF0J4W2EuEgTeX0ze9XdeUpCF2xkBHNP7uV2N3GTlk+KIB4j+7jkhsY2dx97KF980vdJbgsGo4zG
uOJfRMNLmHQXGvGRjv7nzlY/9Jblu4Gtqy4Vj0SehG/gMCmJj0336iNbt7oXmIczCH21W+7dYurA
3TEs6ggf+SurZiMwODC0kXruoyyX0QponZTuhAPlG8srIyOf/14a/TA9pHrB9nb/G0Z5DHKEQNUY
1E78GdmmsJCPdf4ykd0jIgn4XuJq75u07BTHYoQ3ARYsnRPlu0DhdGlSvHnArjT9W8xzY0Zg+Jer
5KEXgwAOqQjWHJcYNnRyFqYgbzHty3OJ+VvcFiC13md+Gk6vWvi1TACP1Jv3gJVzEdWzu9Tn67BQ
qlaANgAGk4gUgHyDv7+OPvmSMW8oSkTNyydV/1PBiSv26vwUMbG8nuoHoo7afI8lb2zMbawYptkk
hTZ0I+34wL86FJULhABOu1P7hb/qTul59vohj0Y0Nua42GbOp6sKLYzK8IYTr3A3MTiQ1L+W7LZZ
ntAA0/XUPpQMSDLrXgGWYEuW0aWLtIurzrxs2DHZStlZV0/xlnwpvGN0ewOIlk/Mon6TOIMsXgcI
EWRb5GSaUsfmzPXal5OUP+XCRqICFC3M9JkEfJDQyndryeDVLkHt51EOT3B53uevoRpLVioBT4Rc
NKuxFqGQ3G0qAzYQHKzll4MjUofY7IGtn8dA2zzGxp8e/BORbyy/CG5fCfEkF19hRHSlT5RcH3d2
DFeLsHodsof1+fJIDMPWJ7jutnIr7hpqmiiNi5X0TVJfVGDdx/dVYPRs7+1DLRXl2AqbGTkJ0vZc
4iwa71aeTcfTOmsKRtzJPFXTrYVGLfodmoTdajatwl6JjfhC8MSkPLMVC44dcR114A/PVXJfbvUj
UrF/H/qS7YuWcca8M7rJWuV52wKDE8aZc/OT8FtMKDNW7XuwswK45qUNKw/ATJSLnMw3+UyWc9/r
QU3m2b5YTYUZSQI1kZ24LvZB6jd27nUV5913HDDiRi7ku+L0+vT5wto3u6iX7JZUDAReX+OSD+pz
fAg+6ypythXSfX/K22hX7lc4aa9zQlgoPnb7UEeTI9taij/09lDb6AtogFNK9e9Fc/UAC0nciTMY
XYPbU2lFx8CyqNwtg3RPK8CqHrqRoASp7TYEirG9rH82pWKBla5Nag0n8FfgWuWQEBF9U5g6bzIT
2BpyJAtbBjBj3DOZlrsVN5xj97zaG6XeYHImRo8fl6WUPjMwjz78Nfwbz3XkBsZ8fsbFQQcBnjl3
KSzy1B96nzjoI/STjtlyPSEIBeGXlRFpySoQJ+DMgw2uXy8V+py+1Ni+qXuMGQcqGo1CZ5Re27pZ
ahHpoqPJ9HVDKaw8GPqHHihUlz+51+zJOhtAJfN2IAcQsSCww0poJE3Y2qgykv7CNTH+vx0DNwLj
WKaJ0Exh/ZREGmJKJnTY5Xyj5FPzcgjCTAfFZanqBD2LDNgfXQsLv9ZQkJGcMI5CjbGFfvUZe0cG
WhpfpRxAYAp9ctNdq1qfNRtK1U5J9zZV81+7BQdLicephb/9hH3qI0EyYV2xb4CuSiE1ViLsomgZ
TiNruXuqmp3vdSoKhxLn5n2sMky7GE1wZKcAyrgGhZKKuVtduDEWdyDXIwIeBEtQ9FxDmNY+9rHp
4DxFnWC+M+T+bE08RyyYBeT4x81CITVxTGycLPS59ef6eKoAyvF7n0djL5ie1ds2aycasrEQpKgB
i7uRlKEj7VUuaMLqSBdYk1GqDVigdhUtIyfcz+PRLxRI5DbEzZTaPTtM8durpzdth88u9LrJrXXO
+K2WjjsOOWF5SJHi3Di6We57EpH6fbRs6sUIdpQtPVg24Fp0PXoVM8w/dhIwcOXDBSD8FX4eGQ2J
1tGwsRNKWaYmwW35N1MqNYxZtS8Prh3wKmUvmUisDVKN1FRfA4G5zSxxrAcT72sV60E5/I6heHTX
BKarSk0aO4pppEdvGhphjk4J+/Y+XY5OJEXhx9snJTrykyagaSnvsjvLL0T6wAn3zHrfDmulQHIV
7fNeeVFLa6cy4cGy3nWDiWgWvBe/byUCeHy1oXJA3sLmwuDqmmRnHOXWM0UjI2FDUt1miI34d47+
6r/0oWvVmGOL6gRw7qOv0JOZoGUBgtYJqtUxR8Zl+HgiEsdvvTTGndCq64t1GLNXYEkLP1SW1hqr
/E1ogRPoPZjVsWiIf4ooTr+hsaaNdDaUkdR5uzK1Iz2y3m3Q/zo5v+gGujUyYCULeHcXKjTUWo2J
FVUvXVQXINllJHlSg4F8AyYnRLRIIf17ILaMdAVO0BCZrI1r0mGTAd8K9mXDnATIpXLzg2CbbgBX
XeR48/wMWrvGME5/nDLGEQB2iAdpr5/D/T0PUJgJl0CuppagrnE3ilh2+1VS5CtA6FIm1DSXFjol
bxYHX/GgMoPJ6VowE3gjqBXZKGV20HGMRkClp/RmW16gr9HdS8VBMefz9gZGEDWiqk6ho2zIZQH4
vD2BCei8x0MLzGg44JRKeaBn1s1puo52yf8wI8ZGHmemLQ7tGm5QjSpKHyAN5CkBHSGoOhpcNxZG
rP+8Pf+RwgFBj09eaPnOI+/M9I/SU9PuloBtEnGgYUZcdNegU1YXav7fIUSG1n48YHdhxTu+TCjf
GL/QJTaKlKtBkEtRZOsfeDMJ2sj86NMAU7xXthwn1o1/nvf3FhqejlYZhIxXjla0VYxP2UEE2SrY
YDBiQLCBljn+mfelwM+1ORMm4MdVi9sYa3m1rXduPKHs/fQ6R9BWLSc3gQQaNQ72iF9qMVD1LLgM
C2F+L3/AenNfrG2p/RXmPe4BP3VhmQ0pryqP383SwgGBDFc7cAS5TOkL//GNPTZ6u5FjKOIvmdPQ
rQzFLZzgPgniSDVkaXDNpCkyjgAnZKAP3/DfPzi14Gest9Agdrn7M9dQQRD9gcqp0RYnLpRELwN0
1B5jCQlreGNmlPvf/eumJGufx7wfqwuOkDQfX0Xtxad4ikv2OiG8zwYEPUGb0FO3vtsP2a2hNMCy
GSQCV7YbGSISu2dy4loKE9VgpjPlqEec2mxp1i1ie+Ys2LA9e8NIWRFM2utboqzcoyNBpsoa9jnb
ezcwOdnpbLJ3ceYZtF8slF8EzcaVGvXqZvkX51MmcHtlidg6UEg66lVijCqLtADp7XHHDwbOqndJ
6xLATjJ+Be0OIe4Mjc/I+BwnKo9IlgeRWcggHEB7j5XvLQVCJ3Ixjc8/lG7hcs/ufG9avj8GIp7q
19qWzSsov7uTQZ+Q+sJ/U3EqguTnw7Cefmltz4M3LvQrr0lAqotUKsW2w7ZZJcBUMjm3FM64iPBS
HxzMK74cRJQeXgLDjguaBnuL7TToPsbz13dIkqTJcgaMp2LBXCRa1f2S5ASF/oc8na+wennIJIGv
ZXIfcon0felxmByAfDETBIRDYx+QHragzzi3Z2deX1fBxnbyjH7NgQKxkUoa0SL9JPfET8iYoXpE
AhxY8NgfCiLwYX49Gk038cjW0xDXvQ96buvnCufewGJJOBNsUKrDLzlWeU1A7Ne9CsUDVAZbd5yw
QaNY3U6Cr5sNhuUARCWnNnaxwMz92zafrsKQdELkcaC4ziJFzi3zasVccUa1MFsUDq9ZHD85depG
5/V0W53Ap3icQ3r5/MUOuCGS3kvNpbpADIHe+RYcRQ0/k1vvYsrIqgSOXC6Q2rkxXD59ZzTqo/QP
NIuSlyqgf5dp93x+ZlT6PXbI8WMyPErLHkat9P0kp3USV9YD8kFiWEjVH2Ot0QLNxtU//L7++kFR
otCCx3L03lN+jmV/cny4KNPwlt2a4SpN5PjwWwUYFdWB7BK3dTLqEzqdvpsuTd4yM0anlPhPOElY
8qZVA9mKGZyZ0Ni291/7x8c49tZ58GOL3MweLWl2LNm1ClHus7hEPkbSKqeogCQAEz5v3cJXQXk1
61M3a+PxCukPoDNpbOkr86USzKBO3gA+xdB1/P4wHlzEMNVHhJaRzR+n6S9niDXShT4TKit4fmgG
esajqKG+k53X8hM3pb8Ndu9XNRxC9CVgNXNFHktDdWVi6v5nBiqduTFDCu6xsPSXNJJM6/W7QKJV
kjdG16WAYqA3lVtpw4ySgLRXY/W+piGLFifeiAP0LfL0HVU6JIZTHklQXWAMe+2124jrwnnM++9A
vkmNnx/tJ18rhv3hWXL+Q+E50fDKtzLRvCuq7J1cYfmz4K/E5tmpSe0+nnTuhHVJwlwFxfYi/uva
ww/3Bn9j4T+z9vz5TK2DTKr9muhah0ZCANm+Ch1xlTejE/XxNdqv7bOjerPzRQLu9QjJl1pWGPdG
obXXAXi2ioWwZF1L7euG3N+Bvjk26M7tHrZWn9Hb6yzTesFlxYnzw2BL6d6x9g0ghnd3spWDjro6
utuVWadJRs31GmlCZSwONFWrVtNksM2krG/OWNFZ0+On0fTVjCBMbxmJ6TL2/jjPkdjdG8wpvo4U
gIRWwMJ89fstEe8NJF4cagjOvuer18A37AYlmU0uEjDD4xL9CpE4QgXaY1tQvDtD4ZzRTH2ib3Sc
HTr4QRZ0tYA6Os8Wp89eNR6bavVk2AR3ehJPtcCsA+rF6BtHP3NvnJdxkqMrkhqo8Co5DzXNCX+c
TBs1HZ5bQXTWoRRVdsaTc5bdaLxkg/vTHyPUvYYZfcojbDX1qyvbpfT6wZZRLvOCjQMu9IwtCNRI
J4oydqlSxR+RXNIhVXZ4S3XLWRX1E0azBRMT0bGvsPz+uHEsQc1AbztbUf7U9YUVe//sTa0dafus
VlUsMSSfas+xyYHHX3edg7yIGkiQh/q939JnFi0fdqVl3CKsh9922tR0/t2dMkrD67xvhAj9Z9/r
U6msU+1Ku3BMkgvcBfvytYGmFusaBHMvGsLBPEpszP+GjABSh6umKl9rITaT5Yc7Fv2fl5pIblOS
CmUuXUE8k+ztOveusDmm9BlmRE/ImvGrWeySJMMykNY9SsZlDVeKKXwcWI0QUkB8kidPhWwip9zy
2JfMb9ddTAR/5BDn/cuA8UtExPEyFJwzEEwNEuoOa97YQR7FxZoFrgVx31axASdeWBJvAOJpUoGv
0VICpI/UrXBWmIqDMBbkPyXaNGtWEEKaQEAYASWQM/SS7i865ZDpMATCnM8z2Matvt8H+FCkEx9H
wMs8g78A/0fYGxDbPHI9TK9EP5GehdOiqdLUdI/KGIqknv1H5ItqLRDWUUAnF3hXqtSnq0T8LmzP
/95NcaZU00WV4EHK6GfTeCwFeT3LUwWbdD2YMvrQJvFcTdWp8CBS2nv20maHhemqaBzOfGznBNkf
2oTtgInWkHxHkk96mJ+mHAt31J0du9uQURr1sE14hcFOuvsnj6S+rEiFuGLauYf0r/V+epzUA7KQ
gNpiTVI5aTGIGIeV08RlVSk0LhUX0B6DCW9K3RA/8mmM8Stn5+aWwqzhjc3OQLZkHgslXc07PCUM
Ikk/+gK+F70mUEhjbYz+oNNBvYrinD7x7gRhNFkmaigdv3gkYhQ6mkqQEhYTtDBClfaXz2vccGZY
OzqubRH2BISaSOOIn1D5XlNwd0P27HRk+mZukkinStAMBu0jLq5Op5yvUO8IA9NNdXFf77wmcW81
L6xr3ZiFIlhurTUfk5C9MHDTUAPF6zj+MbbhpcPOa9z60aVD/tFPMDg3Nw9liGgGNJGh/VXYequP
gTFW3XxjNuSXvcil7oiCdHbiRubV88mACtKSdzgqdNCAkY8Pfka7XjS1pHAKjZV4P5XN47Yi9SUn
AZ36q2k0V0OmF7vmyyVhnximqCpG+IwF4ZetNgoOF/MjMR+o98iCuh1UkHec022ICfS/jMtyi/wL
Wx752nuHlGQG83mhw99V6VDAGAiS2MgjIuWaoik7V/GET0HfUt3CX9+cS8s1IBPt0Z5G8WksTw38
e+EfgJQhSjFgY52t1o0T750R1c/41wmrF3vZ8aV+qK2ep9hkksJbZjZFP9X+/BSVbEJK9Ln1Gs9B
N9LnNZAGOAXY7WyDkp2RV7dY1bAEWFJgINA94pAFBNbkYjtgvKFmpdBvyH/SB4CGacSnzFTDuWBI
i2KMrYZzNMYm2aYPuajh1pRCrs4FSnOT/UZuTYVigfLxC2zEc5f54Ksalqg0Wv7DUaMUOG9XG2K9
stN80W66M590RPM/Q2lPvJf/XF0dP8bHdtYSJpbwfvOZ6Y8GLIPHRir3LsmAp3offOOqtc5zaGBY
BPjPPZx9XdHq6i1B2q0zZjXIJQ5LFQD7pIV5ayErgEuPkqnk7iBb7oFMDw9UocSIs9b1zd+kclsb
VS32kSbQ69IVf97/3ZKjU3OpRqd6SBmg3G4ySXxEa4ySu1D7ndXhP8NhAB2JLSph9zqz7g5vJH/j
8ypky+O4C9IACOJRdaNp70ltiZmriRg7sWlulTV3VYXVTHNlB0Ls1ChCUOY+ST8aHsDH/k54VvqE
oW4QSnFRACElpW490/323Zsjl3/gaBoqqEEsbb4oh2fWH4oG7xXr67Jc1I+yF35ZOEgEzbZftUoJ
8PPNpfl7W4z0VirlhcHJ3wN3Nsa7wYf3efxPD1/9jHuqJ3YgOhimA+xDXNMHnnFtqfGoZ/CvBinY
qCGJtqEyzJxgMHXapGfkKUZfWRT3GxYBd1SUCSJlAXL77hphAUxllYNiWqct8MOyO/39OpxN8usf
J4XjeyYAdyxPOEqIS//VHLYUgMmR8FVjc8DKhAIIxy3gity7pXJI5uxBsN8pyM+NXfbzXdzf56Dk
9tal+7YjfQcJT6SqUHuEcj1X6+LTCajQeYsvczZZMEoepQCwXnJqyH1U+jEoqlhMt1lBK1Pa1aqY
1SJpBtvMKVKoBR44eieD2voPAXK++LSlTNDLXVsLOudYWburEpzxtQvGfvlhspBACHZgpGOGhDcV
3IQ/t6Kig/w0DBz6TYSGF9qddlkjY9vKuahPlR3gUvphdkhx+G+iPeL7AEC4Bj+sQV9QNH5O2hok
FD+2MSKoFN3EtqudDluqSF22Ua8ZHkAG2FEfMAVP3YznjMtKD0uLIP6NpcQOdvSJm6jb/uI5RUxE
WrrElcKrdag1gj8677A8X/9KNlKkIW2lp67loaxp0yqqavFzEKHsuCJQaAQ5BjQHGV2Buc82fA8d
v86PMginC/qWZtw2DPJ9RHyrB1oGMzN2763M2T0eRlgPl4wbikSOEYqWmdYYUEaZlWswuskGKD8B
FAbRUOOZoVgbQd4ObUECUdkiESX84xFae4gCnr0Wgu3RlHEErfx6+uxV4yxlcew2oD/idSdU8BZA
ZT0D5ERNjtiX72sSDt3QTM/6eBkbgwGV/BPZW6OJTOGAvPVSXHKn5kS42Hh/4dFL6/GWGz0bu+2/
pjcYfcD+1k6S4GjQNGZulRIR+lozzaKi5CPusRS7TpfNq1FKLkkis01x844ROEvRMjgKQVjOBFZZ
OrYQoOsbkOw/ZQj+Mfef4Euovu86ZHrEPH+oTuBFd/WY23tbAUMIGeoHq7eOOYPjqQOfdty/QBy9
m6AYLm0M8gkEUIxLnKzjKyErn4ScW8u58lE8LxNX2VaH5EuuGtQJOSDJq9dbL4d5C5Nw5c0Usdp0
/BPJZARuKbA2rMi6vZp7iOURb4xL6vpQtr+MpKA95Mu8+WOXs7S8bWUCxZEJ0O89hkYv9DPGsWoD
QIF74iHzeWgZqoIbl3sgVv0/3rarjAmyFTEsnTXRp+cXRhjmYXTCCcpfHMKzLojC2EUnuuOyiGiW
Z6diAIbscSZcJX5f7ddLK/CWoe1DTF1qzlr9KCiFiqGrS/9mydJKBjPa16ffA01dHTbwA+9ftlwl
YBVhCu50dF4+R65X28UjWT9l7+JAM41pN6kbFBkymHfcenusjvUKs0iD6xB0jjWyOpCqkUHTnrD7
/r6OKr5sGKv6Wk35J50to+AvaoAYBVdVTzJuiertQ6mb92yu26l/kBOAfNiHY06rifQoFb5QR1n0
J/xbi74Ve5oL4dJjmVxvxU1seqTcIv1om+ZW8WcMTu5+SgueXvjXEhzAFA52QUa5NeuBoekb15cX
Ptjnv+xsg7NPhWp/G7DRJCAjKnwyJkQ9c77E/vtztCs0si+FX8b1pzS5lLWs6k1zewWX+Ppx4ypO
4SrTg4ruW4Htz5GSdH0yXtLnyc+dNBwz8PNZo2Y01sBEFc90z8GKJm4C4FjsDjqa3cb9Od84Mz7l
48jFZpGxKryzw6i1E8EYUyB8Yyfqmni2e4Dq2Ae8zKcZRWfnrjA5v8TaS0yxaSr53l9Cc99fJ30k
cjd29oZ3fPKPUcNMNKQ3w1jMOCCny7ADSQPbsmlyNwFBLOG0SEHbfzp0hqX4RADhw2VvhUA2yFqq
y4k0bgSq2+1g0gVMXZJ39dVA/RqBksLgV0j2WFi1o3CX+86AqJi7DUfYPsn2Sr9Et3m9CUSh59As
eM5tQ2jko9W1rJiWW7FfPekJ4mHDd1Kf+LHRq/xxLC9fhnv0Rb9Y/Jd7SZ+rwkNfpzG7u415nIPs
iBECFPkiC28Y0pEDyEw47fNaWQoQS12ruP18PQ+pWoam/rcTVfi/ra3vGD5btxYALQZjYcXpdKyj
d71XKQhUeZxPRxcNGX8gqxIx+VtZIy0dMUm4xSm9LA9cL4GkqNwvkHvWbQ1G6isy+rGKoMluQ6n1
J8TUGypMUaQnHMlYLmp4zncwgq4h+y9VzeokOOdGpCYYKlZugPZQuecqQ/UP9pMroXfJeOv1Y5uI
DXg+TDBXyvEXuHerwItdZ+G1m4G0v60rkahSzZLcQ6qhWk1r4XicWEWQx4uUII9q0ZaZAIekVwwa
mf9d7+H9oHZNrEXX2QRbbW9A9+DkZh0Z6HdW4/r6aMgr37Ys2DTB0AFHj9UsdAvSbrPcK1AQ5dGK
Kj6PdexUUW/vJtrDIbjlEPahyvYOHsZsIU9sk6LLoY15oZXt4/1AVqhn39sJgjbkj+BaaXNXcfdc
NVboN2faw1uaGd2F94UexeupfnOxGXBMwGiEuphabUOSBGvbTtnCmH2qRqmsTeqppzqtNBhvvWEp
cXOB91D9TWS4RtnCObxN1BlxYcOPNlP2Li8yCH/Ch3kr6nrIBBXThCyfx+luXZOj07+vrJv3dyG5
Z+/WptZ/Jds/sBROXgBYH33ji6twFYrY5umSRACwC6p3B3VIhXs9PwVHviHpqnJzjCNswwaU1hDM
k8HyglanDYJ+JTjXCHsTeOellvNOVNq/tMcwnnX94vb7lf9z91m1PMjl69hg40Aj/ex5wdpL2t8Y
/mizkyLmehg2SyQbv0wQXpX//p5+QpUq3jtxEfyYOqTuYye26wvTigBcmQM1MRdllX+ZlIeEXtvs
apChWPIySTqo9Vqot2FS0as1ojaAmC+qPdd++SJLm8zmW8lfm4zVoaxB1pGmTZl26ODCLtmd9i4T
alo6drjCnIwEJdZRrp/VPQMkEvKU7TfE9DsMKUvSjToj9NLX0z7uqti2WAtGmK50W3vZeA9lQa5F
kPlUlqFi3/7V++TWAgrKZnTHgPKrZVWIxlPolaY///5t1OhMwZMV/ro9/cby3UAetn6d6nIRcGOe
8LsksWQwujZb6jGRs2EjGDwIPGUT4U4R7XLZp4KIhutghJBsQy3FAkHusYcTcCCquz90V1xZe+Bq
ETWmhTF6uXLjifTmvF/Mtt1IvQY9dIA+fX3uFJyjgEeZzUd2JA0gLytJcPgriU/olI/OUd/UIWFG
FyzbkKLAWyynVjoU2KVPBqUKVC17lUFtFzjId8YGASBw8IR/0tHk8aUF8ZA2AWCavsC2CcI2ef6l
LawtEynss/u3wHMCCsrVTT9ojuJfd57XygS2aWnV9aCHNDGg97RmFBAHnZFeN/cEMsmxyuIaxtgL
KwdtXRXH/UMIpBaZqudud64WOPgVKvQV46DHM4OWZKRx8b+T4DhLVJ6/qXEHWzXPNIuns3owKQUU
0SpTSA1tWmw2ltNjQ/1ae+ntU7wCv8ujXtfRxRaMQdyBOuob9myLVmHZ7j7z19b3POG8mXCh9vH4
moOOuz2BsT0X3vnQvaheOAYDDgCGWug/jjwXiVTPArCMH4q4/VXKkKJqgilJfGKVNLP4p3Sy+8g+
U7QD9drCw3MXf0W04bD9I8pdDOXImHqn0+p5bkAuAr6GlUw2jFVc6LIkfCTKR4zBWoBXVD2CFp35
Xxh/EV9G2CYWm2IUXs8cLO8VMTOXrFZ/OKaE+ismAdUPqNAxkuNDTuZRQXXOwStrOym7o03d1MYp
IqGk9dCjujCw/U43VpZiI7JDgVXKM4pFFG+R6L023SuZYO/gM1fxsbQiTDCzKrjnAPm/C/OnTDbW
XRe4Oec4onrbpAJOcIKdSCb3XTrqlyjX4bX3ImbW0hXcMp2mHcfMofGerInKRrKhQyyDSze8K7/S
9LUMCTuwBRevMCGon0R6vxu4QfoUx754eGLuFuwrAqOTtP5yb2wfXpDEcbxbIEBbKyH5OhAne24q
fQWjlRKiNpymGEgYEs5yLANGV4c1L62G6hAbu+Mvo/hKkS4NWPwpwDOwITCB9oYUmZJA2gXqxfxN
0C1phAKRnGZVEqJdYQRQ2PID776/V9wpM3amfvtzKegSAB2Q4l8qqOUe0+eqB9fS70BpyhaW2AiJ
lDZONGCJAdBuUy5S5zHs6VEe6vPHTxo25BffblEaC8eo5KH8sY43Jw7pyMkfM4EN2sbp0YCYmXIn
SYi56YwS9xpibrwXhrkO05jvfzLlpABc33Ok4GKjVaTPgCivL6Jm0Cd6XALplw8do+ZuNXF+mpXN
VszWelbgS4G+OppbW+mw3SqXuUMfISr/ErKec5NUarZBc9moKVRI2YDM6yfQKyCUWCSIBxg8CJU8
JaJtGtfTd/V5lrsVi8/Ta5g24d7zl2oXVAoOfHuhXL98622PU2mUgZojR7DX7KdiSUwiQcavWkLI
Umr+h6ANJk7sbGDeg8nnKzPtCi265rmISJIfnYB7sJaks7g6OHg0xPFVH02nU3uUlCF3PcDZHA7z
6JLNqEnLwC4a2v89eTyStQKpTBtD6nBtoNPYYnUkzy7ZYOCUkDHy5SzKJY+CPMAHVKKKUjdAYxrs
hUOmzUiiZ77EDl7ZdJhli6V0OaMePcC7zrM3IajkPTRJuZePMb7Uf5nBE5SxPrSiYSg8X6p7VG+8
cpkBzEbEvYRaVBsODR3ma6upC8FRq9Qzb801Sz9pX31b8De9vpZWPTxDAU0XnwjHenzLsdZ9P0A9
iIIrXzHbtEnQl8hj0WzN82obt6aitXa3CTKHNrlFwtY93ixzic+1ekLLUBpcmRqRCUNEX2cs/RvE
w9AffqjzSZHFQf4TcX00JIT1DAccX9cpi41sqhlCi2c/EMYGpnqJUQ/LnBjfQtG5vyd4+wV0+gCI
xfSNYb42lToHre0xrc/THKsLIEEVHYGYcZRbqD54/YClNqKduSVA5JZb/kzcNZlsfC427uNmaFwb
B2xjeo7/GTZk2saFsKb5j0uj25qEfqcY/7uECskWybPY7Rr517zqCYgw6OJYhJCJtf5nmsv81s0E
GCECZ7gYppdcWxsn1uZAHLrzQJuqnEKoQsSRwWuBTQz3zJyNeqiPVoAQ7znC4wXZxEnTbeckCq1o
k0gxNxzdg0D2UK810QhCr/WHkx5SEZBhy1eDCE73IUQV+tGdcYI9hKEgmKpGZOYyW3iQL8N+zMdn
HBrLOfqkCUdOKleNUHHg3eo1mddZv7fYkQCueZ3rx1w5LPGulw8gIq981185o5PzAhp3JhBxx6aq
gIF0SPS/dU3fK9URogYVsA0nL7welmG0De5pSCCJIFD3lZ6mmUYJGlIcAYFiyUOc5FG/3T08tHQi
+y0p1SLL24h+noqbVmOsfp7mzQHjwflQAoaxUK7UOxKQ+KPKrl/L9GF/MyPqIZtJFgawZoCIrQCT
JPHOHut3gwUwpG5Twt+x0kpu7djc5fXbFn1YKU4zTePnjb2sFKP5quJdGynC/WZ5xxFsKO5xN656
ItL6eZMfx763MpE6ZW1bo6HOoUbrKS7pudmXHN4ZuQZ2GitxoxSILcvGlSZOgHivWMxiY8pJiYpQ
26n7MCSGIr7jVwRwuHg8T3kW4+EYwpRnzEnNXUyKYR6CgpNEqdL3I/o5oat2RqrQzlNegtQaTAf1
jj74BJAjREqZR76UgWxdbkcUDUNp+/fj+uXRRDDCd0LV1hhHGV/+d7KVb4cDd6IbGbavE7IZhuIk
xQiN0r4pSVCkG5GJrJuugaULZqETMU1i6ykgIX7VRDVTd0kcfaqS0uYIlXza/yArtqRincsm5W4t
Na1i6l/4VUPj+uCekuitnDdb5n84mM6rAcLmq/0d1IOTX9JDJHZdM9N32kUTraEhnLk8DJNJ70Pv
Z4I/0FFsRLyC1m7YFknsVx/JKvo1WbB93vMxs5vI3iP/AbIqBuG6lJ5/RIkFzQYjJ6qD7UXbVjBt
Cq+PEpjIa6wusptPTBbr5WrmuJFtLD2KjafsemPOeRTNmhvzFxnFaVMPtQCKrIT1tHYqdON9TPrR
OohBw95cRD8k2Ni92Cn2m5/XmHZNESQqlQCGsVqV6FrHoHrvc+AJJW5hw0QY0uG8rL44hfjYzUi1
gsbg+56wIFBu5nrcG1Rsb3M/i0Wgzp+RI+k2mUk6y4zlsGyZJOTEZO9VAdACzPHDejctV5MjRfQq
GXRemwKGAyDlqTOrsf9w3pn85TtsXO8lsIqX6PyJy+Eu0yn2uPAB4M9hJYTs4twOdgiBrwlKr9fo
830ILmiYzwTxjyA0h7q7k78fm0g5eMeKAukB1CT86S2UeDWQoR7MamDBGzQXLJkefJhYxr186vVL
FOIUPEXSjh+hD973Ah3YSOvZzoV6EG0HbKbUirqpReGcQJqMA5hPcO30BA2vn2alMSAGjrH5ci0N
ocVso9KznostpNJmzKUdVMVBCww7t2vzD20JI6nT2WUblsKAaQMwQd/O6L2KuWzOiJlUXg4DYTz9
wBTZOECmQA8N/FRTSgVtc03vACaC7uvFA7/UcLaiB3dLuviYA1A2v1CXjzHIoIzs/K+aZ7KFgGR/
OMyj5oDybeztoYOViN4/LYvl4b9o3fSU7ojusVeKiIblYffi2b2nPwzxaCi9/hSPdbE3rr3j/bjo
dosiyQ9v4D/M2D81xc77cscQCE9KuVy9KftWjaxyY2Zu4EpyhMwvDDsOqg2cLXpsCGeDOCNHMVGl
W66/91El9C9wAgoD2xuj2ZbEVH0GskgK7+dXZtgf7VxQkKZNTuDCvFSn/d9ltEJes8vmq0LOznYO
GJBIiD22oftXGZDnSCmeCLwwc236ySeo1AL+ptKFagoTj2AZ+uwDJzThiUvZx9kOssWlw3CoVB51
ir+OeMk6msZi02B/zupP+F0cHjWQ7ko3ocGmZeOi2Iw7ABtb3aLC+v2PMLbW8foQj65rUcbZOkOF
fKPoSeY33hBRiDxUYiMuoku+F6kx0I8R992YGAEC0DENCsqXXsqJ0fxDG6LiYBp9MzhhYLoyN3Y0
FkArrdW6SslIa+dlOwD0l2PBXegsqj56yLcuyloBeTmbCRMicr8OlQKHeT8gvtoDeh5riKuGBRAj
o3Mc+appOJKClNjMPQE3YQGFXe6lV0FrtFxLo8sxnmzxk8QWNl8QWsl1232er4f6c3XeaBGlUj3f
eCfD39lXIe1ClwnMaIPxnsI2YSAeIEt/3X6vpx78FFjd+m1ME5S4PumdrtIpHR5RI0M7MRHLUZLm
qFyXFdoNB878tfCotutw8N3FyEiHTIEqwZOsyjgIc1AvvZPo0odBJr6ldOCaQhBMhzqMnfU5NNGU
MFFryyjnk6Gcbhoc8G0iC4qHCeK7rS+ok93c+5yPzPnnpnRw7aCBYLfPZRFSg7u4bXKPX548N5DG
gupUkiyhZAoYv3pDEvptqVrojPSKW0YFNzWzRJaKI3k+Jy9/KqBIwphnwcJVAqRNlDPS/CFeQ7xI
4zugdacxqLDIKxlU6lT6r82QEfQ40JaQbGEAR9Byf2DHcYbVPifoES9jNtqK+7mMsf9jcd/rrW+4
9/QMR1njLTe9cTwnIl+zm++GaVhdCUd1G9JDsHGa4xxDh4fdokc3pF0VYFLx3OhPkUQLs42/OWFt
VCZhNoNTIhg/We8Wf+kVGgVWt8RYxrk29CKfxWjtseOEGYouE9WpSN43+KZPL6D6+hdyQbdL8Zrq
OdGan63hZJnuj6mFnatvIWNucMY+mIR2S2vebma3lHvLUa0nKstsyJ2rp1tGg0mKu8EuyvprAfcw
vql1MbYKP2ZxnkTf8598jaxQDtzENcTWIe566lwYYU/LtdOXWGz73AxMA4iZvtn5QTYmyuwIn5DA
8ZDPUqkTzRI+90XdYcTOI0N7f+/tmOorbmmHKUQ/m7hNJgAALP2XjUYX/42PCgA+fVR0D6XLH/u4
Tl1l6uFdWqo9J7a77ZXYb9evp5ad7oS3bUOHpPYWovZzeK43xG5WM/YrokiVMsAGjTTouD2NwqBj
9eD3ldRly8uYTonvlsHwCfy5jpUkE3QRpcd3Vk+C6Y5mtb64eoG3c7cdfQDZjjJ1VydZw4SMppNj
RufkRgsGPVU4jBhkhnSU773kieHwinFEu6ufEGzHy2wXG6hVeBz8qNrCEEb1J1ZgK1OALkR4JmkS
qDmOuxWDrzEy6jHuZ/MG6Gcw5nt9iFlCF1S83UBpziXqDwqZDYDSuaViglxAHEak0dTF9IRTHL8A
zDMeJqga7z2NzQo36+m2QdbykCoF3tRce0CDQiSy438QQCl9ke1zZ2Ob3elftcuivkGC2W/nOhQS
qR2qVICUeDNEWbczl6FtQ0rIvGI8wWeL7DLKgHE2CHEUdWv31w0RDWwIIY3pkghfZqGPeuaATvZm
w0yGFEcpUug7uQpc358mPRW04H/Z5Unn+g8H1cucLh49CMsYtGUj456m5oR8K2M4E4pjVZKElcIf
b4crZm2jIvceu+94RztVbFM6LAnmbg8JOeVKg4BjnN98vrw6p8rpQjMZJqL0ZjlaHVZoNd8qo6nj
aM0huS9BfYVm3g4Z+tNH9IGbtDWEMXV4dGFTiBwgjIPdSzAg1rD2lG6t2o7wvvONaHNgT7DFmdC5
dSRIT3rS5cfg4T33IMZ1+Iw8LQxCZEefa83FMWzDZp1qelLaTQDvRiA6JTYGsS7tBRSILfOdSJXG
9jVO/BAiJzOl1+CY5WKj6LHf1cpVWM8TutKW7PxaxIM7ERYpvn9jtZiCXV+nNt8Bws8N5UocKkIx
AUqvcCFRE+DtbY0B4k7BITBVAqtvVhUvG1rcU5Y+WXoDsAWlK5mjuBUcakejfC+HkFEgtQ1/kF2p
ggOgvQLDY8MSLYVYYcWd3GRTHfN0FMxzcic4cxvJricmYZ7z7m6kFS/RsWWkHpocVNNEH0Wbsrwi
1PyZEs+98SAsUw3GXFMR2Rt0fqrbDH7tB6xHISZyRAgiY34T+zpncCnPRYAQQ13JwEpGarkoOzYm
K2Sx2JqnGie3UpBUd5oXtOWxl+B3xLUsUzMHdqIWxODZ9sI9MlWgkx3EM539FZjbzm9Cx7thOQih
VRcZpnoiqhsIID7NWf01o+d4mY53JbRIu6hXqd5CUsQH/v31thl059nWji03/F4WXckYRekuDZXp
/EFk2HeKJCa+RyGWTEqw/VjoaEo8yBSuOT0PWgAOi1P34GnyJRAgf1aoJbuwOXeKsuJ11OiDxaNP
Ia+TtX/pjR0yosb/T9lGL8c23SzjTw4pAj/Z2a+3/fG01Nb5ZbujUHANn3vmSJX9iaUjX4HXxco7
C0i1Orxx3SJ8aVng2vdfxLBWVSIRP5zsTdD65Hev2h1DwjZVfE0+hFV1bsxbCXOlGCFGY8Rmtelw
ZhwN1dzmc6v1Zlw+drJYG1HIo1xYsj3g9XuVdILwTS5XYy9ZYFxjxFbBk7/ZP3kcmrpEvlqemIyW
wxklmuMiU/Zv3S/SrUmCggHCFNTItRfF7seks7yDQJzFUIm1B4BCKS+pFCaIO/TFrBQrP6hj+eim
ygKXwKE0Zc1Ps0dKND7m3Mioz9cQOtnV+9fCOIvdXdMq4Bd+JpUa5ozRRH0XgfwP8xrVKqbprMEf
Vg61T2g8qVTwiM9gB3ccQzK2371Dk5dCBP9e7ijCneT0iZKNhX4vpp30Q2zdnr/0kkEyI9WM29EJ
UF0Z6ZeLy0cqH7A+Q9z0TXdRRsDlQ5bc6osGnwsabt4xcQI/SQW6ovMG9TEaPXSya6fFICTCPpyD
7f/KarE0f2fqhb5z4JPtulC4i7CtArHTZB87THU/nUMI7szjG0HJmcMfGuah/ga0kUXCNvMzN/Zi
Xwq5cClyrNCvr72ayK9nmtTAXsxv7jbqIy9eLF7u77uSdVmlThGdUN2xU6Jnvsqb/3w+To2YZHfd
MSZo9gCrbT5FCNS5WSFd3L7HvM6iE/3DNJPYn09xvBkBWqOfAJMdqTd2tfkLGW8hJVP4XbndLnpn
+gvDxH4Ae2pbnfC6QgXpGgZ7OFl4pfRjChPp2CkiW9kooIm0Kit1otl3FGR1z8lGzD2AbfeIZuLo
NV69qRjE8iLJB7yQzqTm0U35nFUm3TTkHj/fm8xnVhMsMECAa01RZb5h+evPHkE7HmnJLKAceIXM
g9+b6vlDX6yXEziGk5XbJm3T3kEEtVgnShruOCrsU2TVcynaWI85UmqXorscpykm6Xna5ijOM4JK
ZAMnXzN95J3etj9t3tBqceQL0bvmE0uLkS2HLMYSGSKvmgchYlG7PKBdYoC7qk6loJkU6MBmrTNg
xm98Y4Ty4jsoJaTXQzK2A90d62fAPU/MzAeh6Uu+yXmfEKS3/PAi7mAbZ7IhkbWg5Db/2F3aMcT8
sqkdsFGOwcAk0X1PxTTKpT4lHz/omc9xUZTsJOmYAKSD0HhTgiNebbsmJ8dY8M8QymYKC7zv6254
V3VYP7PzgzCX8S2hNi9FLgmm8KigZUEKx68AC3WDCskQ1bAP0KDoG39IL7uSg2m8YqCty8mFQ6Ps
mhoNND4Ex/83c25t8XiP5OTPWKQVrVpG1t7TOvFgNApB4QHLLJcAxszEzkZfSqiKmJ6tvzjRILDk
SBYlvyEm7Bzv1W2NyWOw2A5XO4EQ2xFbksO9yGxnGJEdtMQfJRSnjg/u0Afe8xOXv4WWdVV7PfVO
+KtPzS2EcqVTVGyVIOPLMnwvT5rWN5hLD1YpRHM1dLW7KMrTZ50XEdjLndGx6Q/G7OOTu853otAc
krXTjYxvj+1p1mFIgTqSiVyEc5fDbj6wlBmOa9XgHQG44cyg4ZUobYFMfWdbLyu6tMugvsm4659L
3Plz4DkqlUimL1Sr/g8Wv8LXWy8hRwOuAsd6GaBdngr4KtCkxfZYwCtn9W7J51EEvrjjeJEURqP0
kDHKPHKy7idxr/vAcYfoIiElqLj+xy4I3hjfSNmXmW5q8IP+gvYEWJ37Vo6oODo1TRbd/7r9BYlf
mWsjZQ9fXAy/tq4bJlBgzqa5cgkqZqgB436pKUWLGN7AKPD4LbT586yqH51OWx5u/G8GoGX9av9s
9ti3UEkurM7M6l4xInm/gMq9rfQ1FoIho2VlnE5s5W62pSVrHBEOI4m6dDDy23nAz1xpKu5lvDX5
eRYMV8fN0zVGFWHZNdl9lKTffA7MeUj82LlJfMhM2RX61Jz2Il6WZ3SQlR16U3i7fdDKlAU8V04T
bUIYGiGxsez/fsYGsSVi7S2jjISwvqKnvdQaGI+ZiGsaw/g1HHt5EtpMK+1UhrbXdNvYHNky8uux
k4RJExo8SanEGOWN/T9q/Wl0WNbw1YKyjNrENlfxwiEnIqmX9nuKoh+Cy22PlRG7o6DBkTeXoO+l
OfFAlytFpbb1ftGPqohmt117gBme1S7Ow085Io50/SXpJzoP7lAYpzZGe8Mn5DbPM9d34r6AyOak
qvKo6o0A1yz4KQ4VnjyZ+6c5cPFQ7mxBMfZGszyto8mPnbqrS+j2EEYdacpbMzblm7q/8MVkMB3h
Oiod7+OabqmEcHfrvZWEwx7J/btq7cDwb9o1wl1a3Rqw13pF6xr4PVHjIaWnfvjb86tUjZTYW3nG
ElRAc18YKzbOYRX4rEGIeM+B15f/xLEjJVmAooUPjDdRQoGaHapMR7425m4/TzigB4EEZda8Mkcf
d4ZIQEfyTkV3d1MJi6ZNsAuX4gXI+5lbf7RZ2j7Ff7DHPizM5xbmQiJwJ/dgFL+hQa/vmp0ISTdG
9XfoZPFD9pZI1ScZ4Kq3vu7CWQlUKQc1lyqR3iyrV5A5qd5+Ftl23pdpXQ5CM08yzn42AlTaL9VX
KMJJrXaXCKrx6abgxROpStM905GZpdfgtVqj4zMEqyYAhkeCSQtFxds2jBL0b00YRN5GuHVhXoJx
7GJIyZBVSBAt4ABoteYxRDs24jZra2DV5isZmAksaZLyh9tf+P31shKcalKnHIZk7qUvmSeOqlwn
eOdEaeeXBfjGj8O3Yj6kBfbM5SF4cqkYFzky0f3RNRIJbE5KGpVXyfxCiI3UrSCYhdgq3DAlQBZy
h/sAeqk3SoDYgF40knIbN6QysnsgKoZByvz0Ko/DRXOMaFzI1DrcW1quPvbGoTNPW87BLRnRtJ3R
kGscRiX2SrxmfHrnljfO2+lRLABsgohk2xtlt6hIyVVoaMnRXO8MoSPsmaNOGvnHwfyXBBrierA5
hNNlMOLDge4FdFm52UKU5SQcLlsrCnTvxfxAucsARpBP13+OgahlaVP7DE2BGvApKT0SbvF4CSJR
f0uxQZAD4/vT/yO83lY8tlAvFQ7Ha7/YE0/9sxWIHKnPymV1FZ8D9Xemwm+P1PwisXQFayhqQv+e
nBaOR62HOZRLYgK+bSXkFo7qPDehxsSteOM1vNgjHq1iTMIfUX+HQgBx+tgmLNGvJfvsFS9YXxO0
vo2VNSpT2SHAUzWr+MOegMzJBNdTc7SYFCFHxng6s1F3zMZR2yJbtZ7xZ9oEmXs+gJpdnDqtDWHF
+pQXHIbOrXcB3GPYIgrS5hP125OR89jNy0sh/waZvr7kkIYX4AmbvHI5ZjfDcmpyrKnkwcY4Oehq
vl26gJxE9/4zPHJOwOBc8r1ChUdZjDEsu9LpKkda8ALrLzR50F73yuWu8P7ujQntF8nm6sEUMm9t
icdPD0N2rad5Bv+Cn/t4iIoMvsgn5fPWsDhbUnEuC9bDhtR0TsvtKChhOASOwNKK6p3IjYs9Pi48
H1L1tkyR/BVHpqEY/XlAM4jTRrYHfN50oAPyJQFq9EA/xdtPHjlbT3e8wit9nHL3c3XalIs8MWFY
shuIj/zs8mQ0IqdY7RQpEzgsFNKoyf1NNjcoLOfYvEWDgIN4O0IqMCKrPLeglE6ZU6zzK0vghyxa
lwANhIHXz8RmIga/4s9zXr96oXvgOeKI7QKzL2KnFt+FsqNUR91C+Hju7f1hnLbm/YWZx/P0tEO0
YJV5jEHE08/qEnTM6SJDk2HOH0YAo+EmkFO7bcMy3HSbzt7vP7dtHyg2wm/8400Oc/oYykuQdCnG
/FhrZT4cj8QxCKgaj2La2VC8EhtsZKyDUaOpfuCTh5FoNkAx5h4sH/Pnt1bEe+uKNuH2kxKiIKSA
Eudje0PUFR9YN2eVyK3IYyVZfDa6+7JdRq8RF9Dk0CvnF5eLLgU8/AsEcgeth0KrRCPJa4BgxDfA
mY2MucHJDb0buJVj8ursftfy9XDHEeg//SBlUgRUR8hbaDJch+o+qH+oqS2/165FeULcPOwK06Oj
pzr+S3nPWv4OCgQSdb36lyZazGbanKuqQIVHsgIMZK0vNPr3qGxONQSKjEvlQhkXzVv4N3hOriaC
vFgVELGG26nwM42Tv1xdccc0cjaNW4PXsxj85Vp4h15oDjSBjEju4re/qMK2Zu1JjnIbV4Zgw+ph
XxZLIIoI3Ndpq4/JkJuhEfRRcQZpcg6Iw1tdGkjMAsVJi1n8SjaCdecMfWJuGz7ifN5X6sea7BE6
1fNga+/c2luM3w/lsQYcxsHURC9QiM/9+84qHGuxfX/pN7IB4xxYmICF0YGjzbiG3tkm+bZZDSB+
Bfnzh4/4K9zsCNB7vHvo8/76SC+xV2IczB9WINtF1pOjLOrTSnjAIfdkujk0YsldAbLVY+vbC1qt
7sD4AYoj/fz9CNBCankB7De//87pKYzazoFDLNaaKbbrAEqA4Mk5jyEBBfrRqKiPmjDWdJMA/Omd
MR77f/OCMcZd0xIZY/B+34OpLoXR3I5Yr7w/Mh44pYT+jK8gDv7qcpR3urrUQlKxG8kKyXv3nHer
U2zjWtLORv6fHPyws7eYv+e9oppD0MrTYtV7vJyF3i9RaLFubDNpR/3xmuOFVbtnh6xevW1t3By+
Mpoa8wKKJNaSCfwIDAMis2UnRvQb2iwvuTi3mmernnZtb0c00s3ogDo1EG6wq1D/zp8j437RXwOI
jb7PcG0bAcwQkP3WIwA88zywWj2KQrvaFBsKF0dGTrTXrdnDf/Y/V49Qf2jZdi7huQHgtYCPzg63
VKKqbtGPGC5idyHKylW0jQaFf6HHtN9m8lXAESi6TvBp+IfXrY8FuPsbmeCU58JEXPJv2bQ05QKl
uC6wTuY/VX0TVHYUt64QpqRe6JoVWqw1zxkXDzZ+cqi/BrCyeECQW4LLmhIQRfXaLC1BNa1ptsgR
kB69cYYEWoPNVEGzFC7P++tUNDq3b3JlAtQR+8IhqHXj7c+glvkuK91NKO25IfXVcNb9WW6QH3Mn
bkAiJBcnjKMthxTjACF4AZNLdYJYtO4kUwXsbpGhhcpnNZmV/frHNUcekdPX7gjVDkkqt+x6lA5M
hMFVi15kDVKfBWnuUdXnG5BuBRxSc5NbBY34yMZIoNNxALzGiZ/Ihr4a3OgOalp3mIwDOJO9trfD
CWA+pInsskCLSmcS12Pn+HLb1Da9JgXsbGQF2p05FfIccX1xHIrY/cAq2KqSo2H8bj4AE53dhrTJ
ewluzTBxxXpCy7LoIjw7TPSzI70c8NDIQFSt3SVAt5ATFmID2z5/dsCSu2zGecgmRQbaJgEiCv0O
up/Y9la/YQaVc/v22iiytRZd6hWDrIbicFUlQRC5WTFMBIMkzMSzAhMAOulziN1pWXA3WuiPEyjb
vvgd8W04fdvOeSBML3eRT19zghq2nLRc1BKeJog0ZsH9WBwxHpa/bfEY+oI27Sa7fVID0aRWX5DX
5yIXJgELF94w0fFI/xen5Y/ZSw3FdU0QVQP00lXVHIbU3WbDry5e3ggCTV/b4Dy+s6+dpDNhc+7x
Zx9Ns+HV6TyAMXaHe88lYPrJSadNowr1p4uTdlVCfQHnAJl762G4mit8b9kOnAN6CuyQQ6YlOZUl
3LEo8ANtgQNk4J3ITTwqug4YmqjH2B1sWw6iJTZD3EyUIbV87JnYZZqTARjmAztz1hezky5OQrfd
OFWqtK8xM1TsQ/JKZ48U9lbdo3vtUhIPDQ03xwTEOJgXl84+NAOQbNlycYK7xv9QSNV1sirpRPOz
cXXsLvVa+Ez/IcPgnB8NS9eitDEXuYqqZe5aq2ejuawlpp/qWG+/X09PG1t9oTD2VXsJVZXS29c4
jLMaX9UGYqaZQc1CEk6ITKMb2+BnsekB2bVXjYcrFWKLX/+8TU3o3RKwiv49ueZpiTWDZ6XCJyCv
/QQvAZ4GqL33jZAIC/18dx2oz031oI2HhJTKGUxc7YpVX96mIQQlwmJFnf1HM82FRDPrJ2VZQ/Un
EYtqIDM2ewovNbKM0uw+MBBdniuqS/4FabLKB1f9igLndXhzcXVRv0/wybxtLk60I943c78s6a6g
BybPoblNlQIW2hvdGsVDEGCF63IsL8siCW7CjjamCUZcbCh0pnLz7cX1hJit4qF+FCTS9nfnvsFY
9nU8gWss2vcn5FFHVt64a7WdZ+ou556GACLQZGqKhw4VF6aJswt77GXT8O78LnWaGBAQOh6mxNF0
qglB8u3SmFcf5abdYrkZtPuzb3FvurxYljgLKJeMh7OL3FDp1tDpQV6q23nKclDpe8BqdHYBviMB
tJdGRkqqDwWyLdREPc99e7zF3RBH1A0XjdeOTvcmA6olEn/oqNbJ613dsu/VJE0XFaKJrtXm7En/
C7+lg8ptF9OUq498C/LRyTjKjsKGGR4CZj717ApzF9U++CUPZN6CbUF2LEgE6YcEVoXMONHQ5rXR
R7BXEXTx03GugCdNXccFH9za+Y0zehb4R9KlxU3K4udNcJJKgDynlZOZGsVjTKr1Mc0wESr2b1uE
AC/iV2vC9T5pT9vk9eaEJHAHCOPgRKeaoRpeu5n1NNufiox6ROCGhneCFqJQc5OIG4AtHwrlc7GO
p3SgoYm6e6SkGc1r7KDJTNFVwTRTt2tQC/J/Ok/9gce+d8x3yTsIm7d0avk9xecZUWI0nO7K19dM
pb5q7LDDLGh5V5ZWLeCMPWgxgwoLUDvPk5vNNo+ugoDeksr7U5SqHZekJWlE696OpAXqptkdmOiO
4O38/xT7i0MVNDkFTppkuR4/oZk2c31AVkxGDqNH3oJdkajYWRFVOyUnR4fkvbIYN5YZdd7Po3LM
XMFeSuvURY9DvKFcpnIknzTkYXqwfRtF3ZmkBHDisvAhSRpOworxdOv7oKncsRJMvrraDhV9dPYp
l5L1UZqXKvzCNIbA1i7j4u8fpJEWE1hvU59cvlOyj0uU7CTORJrRPF8ThCR8ut60pJoU3usp0sPI
Y4UcqfFpRV212mO+z8OIHj+uwa/aEFapXZibosoMc8dovB992YexRW0E9g60+cTc9l15m+dbOAhV
F+AiRJuC9yhDZRMC/sGehe3I28ReiqAuEC0q4c0wMV5aUFNEfFigQRNRjZna4P45Dd5lDyBPH2r2
1pscImcVuSzdvBsBhgObQmBc7PvWFZ57cPQILLf0N00mfNmzfmZADPsXGSw/6KNw60P853zUithK
AiQfloHgGlzSZEEhZAai75NB7mvpbOqozo4wSMbDq3lnB1YfwkKIMPXW+Yr04BzlKjcCW6TNygJc
uI2iryp1RMZkQ5XmK7tIWHhhgRUHXq16aDTC3OAIJzaDDTwGqYv0iEFtv7cLvwQ47nR4kYcAGt5J
8boBhQGfAA3pLjEQWdj7eSDRd+MUUSgeeezdjPKgxTmMd3XNdkaKHzgvhx504/rrLyr+PXUIXgXX
kp8/aGH+ODnR7iEj2aItfeyZYz9SrR9B5ngV4vUexoERRgFmiUrfs/aK9u1bacWZBRkCjafv6La+
+A9tNdG4bzxhJT3mPeu6PlQBFN4fR3h3nAA8FdyWMMU2507BQq6pSbimdH/7kGSq4MLQnDejksjm
d79008CY1KlcnuHzgZyyzb8JkIPBrdVjb7pN6kRBrjrWOtszH+LyOu9V2+nwcxjFXCJf62c13+MT
tlGcBMpuFEdtInR+gGaj+BvxirDSNww8IGCBNKHKFeFW9Hc0Y5YcHLjmBcpxnDepoC9DQfWN2Y5V
wJI0AH9Aq0IeX9JCb3WAig1g5BM9O3EyvMCwzriqXi7NkXNzxpFzzu0jMMPWQNJ2u5DtjswN5ZEe
HIwEK/C607q4OST/0T7ftlKYHn2cuztpphcw3o9hHZc4FznGiG47aR6C4hhbo31S0XdYLIRjhkgj
u6RJ+m1F2caK29tmP/66HRHg0MWeVFFHWayni7vnOIrqIvQohCIo5quKH7sSA7Un4V/FNH1osi7m
/J3wbTkTSavXSRpfzVuhH+JkRp+mGZQAzO1U7b4vkgKmxxX1lG0GiNpq8s3st9pjmggpwOZKW9B9
HKsbcSbdy7r02JD4WkUYKuaCbGLql7qG40LNQ0DLUqM9ynbA6qRd7/b0wA0e0CmmGFQ9tegYqqKy
oO1fhRJAi+krs44FPvWZFuIlwQRr1LTZso2GcACxgS17DD0Rz/b9BuSjfNM/eN/5L09GqzKc09Xr
acJmpMKTjhI2DnN5MxhbTGLaIpCdkyB7zv6+fZzNI65dmhK1xHC8jOOauRR6Izmsc8hdBiogJCwG
VE+EhngKFjwRRuZ39Vu7tJLoC3nn5gghor0TDNdkwWdjsuqm3w0AkEpJf+eX6rEUaoFUvDwLEMBB
6283ym1S6s0dRkwp4YOfwR4HSLYu9ieP8aVQAzr/kRUJkxFm1itbBUZxDq4QiPMvOU5Tffl0oqZz
V+2SAp9+qtXiubtSXuaRAo8b/BcFk0gHYtpBUcGVO7UGg6NA9QiC5WLOQPTwuxGCso1tX/9aBVqS
+QeEwcdKz9w702WyjDMSQH4xmEBLLo1OedZIVQMt1x4Ju1oL01i4KW4ZgDiG8zrtq6t9DkTi0TLr
ojgv5+WKmjzGJPdnjGpCnnKp5TICo7V+W7jWaWcJWlocD4P+72iXW4FV5th0ywCtd2uUA60fVhVJ
/Sn8W7AevzAGIf8AefuEe42vjOs4my3z83AxRCkr9mf8g2BmLFaQYTj5YdxxgRLYQ3nvfaPgqIDq
VhbQ8nVspUPNcm4Hxcm6dpuGsXY5gTyI5U2GBL0YYOhLmni2fAcO2xB5GjtF/xrQJb46/xTAzEo9
PCuSD5bs67trhLxoL0zezrJ9BbL/JSgNXDIPMxG+8OAElK5BTMQn5lE+c0JfIJDM75HDK0Tn8A00
IpIYcFhN9PPhISrrqew4Tian+NlFjyYncJIrJhkw/gMk0T78tg0DYkVdPxOUmfk/NfPKbHtSpVYu
baYVEgr6sWRuxDT+uKpms0uLrYYiEcObDRVVi7HwGUQDrIOLnhe+r0oJR7488F2oYB+psUoJYtg4
Q5pbRkBO6x9yzZmB3EZ3nwoaCIRJ7/90GVuCs5oretMpBxBeGhopD8mjXLILGqztqbJz2LBxAL8Y
KGH+nOeZShy3sfaY0GIUQf2+pGUti6dHLsitwz2MOpfmFrxlCwMT8jhMW+jSMd5uaOShx1y2NKG2
VErXmQg+514+F2GKDORmRHl883RnlCSn3g4OJQDyiEQo+Q+ePUjTK3SuGmr9fMg7IGeJ6ls37Umq
ymoxz1RcBrORBLlMRI556w3E3vatlOLO4kZDoPOq4eJcAzHBcRkHf/XfWR1fon27oZNkFS96WjGd
msp/7Do7ORtHq4SJ0nFsEHzlCSehrlsE9zKoGTYa77EiD9P5m+YWEQvEmj2BlTB6ycQN6wphlVcz
MLfTsc5JNR8knIcLYF9uNBTneCFXyrYGeCcS1dPsmUsxSCixKJjSY7FA0OvzRXZFxhej+ZHnnVdP
hQMVxUqzwxHQ/m1Rv+kK9GlY69QwzBlXNWEtiCxm7gA9raVkhyEIdgLcd6weyd7sX8iyMJBpusNU
zyj9lfOArtnjwD3AhLq8xxyR22jAWnN9MJ0mhyBNEGByv4xJ1NZzhTbmi3PkDdrRPai3U3FdPjAR
XPsbMYr64anfWvTlre5iYKSWLxEHeQrpruvAwPDIcuPkj1aJ5Hq4niF508nYKOm8CUV8Gc1e/0yN
Roca5xpv3B7VvNOLIzvyVlANiBNqL8WzYp8K/CQHFNLSp8ffhMG3rxvBCi2JLRZ4F0mXq1UOBlTy
JrFDPaXDgBMr6BHrBrGsEV4RcVXbs+7hnI6FFEn5eypRqmBxhE6U0PFxW87weF7rxYWbpsyCDSDo
egtOu5zdJ3N/dEII8b+3cJCf8HBTb3oWzCYZnG5hG+iOo2FeWVoXfFGinZRdo3kKSl/WdLyBRX3M
P9I435X81gTcaXOfXOj+6qnpQ9IWFbokvAIol2Wul7IXLGGbQjBELdTRzYLkIt/AQ8AmjrpEtBAa
m62rXuGi6LmFPpyd0nD0vNcWsI+BOrJrBuVgdDx9NVSn/3WTJP9Bl8EkCS5yrwgOq2IYIfaRgjlM
Enh0ML2xrIZAewEqT60qVCpNwOJIfIBIs3nzAuQID/2YoKz663ZZImKB95gKImHZe+Mn55tmkVSs
nDVldAyZDXHENwTFDbosa8ic1FgM2LVbaEALD8yGj3On3fYlCikpSyvwJ5AMYmfhkKn9yzilZfnH
3LJvpj8jHw60oRZJ3ApiMKoNUlrmxah7/b1pqKB/MqJWTB1MV0W5EVRruFV4jYHnxlIEVjO26X9N
KAcKrkE2c7b7XzACvFGeyLYQAe4BpJ+RDPi1MUMzoA7kjlix7ouxeFNuN2tsRnMrBwwZOhplVnZa
gBpJdYYG5wjHPZGrhdp+m+8JAhL3ELvy7jjqdwjmd7oNZqcNZgIVT8QitIpR0SGWeKYkt8/zQMjQ
sgY6AnoG8yxvvtvKwRF2d4J1yKoFtMBpsbEEYlR1YVL7ypJ5kvXohfUMDFWnEDMESqzmGbQLS4hz
Wt/0K/ct17R3o7uaN9yk1+f+jP6NFWJtsu71Pcit+RFdFCEnGClYFBUMWgqybqqS92ms/rLCBLn1
0NXcVTCBC16FFIia8gzths0YvGmKwVf9CAQ9F7nhgwHbmbrNLRJ4BpJBW3LExu/EzPRiGuS5U2kJ
TGBZ3cAhClPxZVg9PE4+73sdQPF+sSjZ/Lrgg2ZcQDScQ4Tj6MdYn63oaxubgUoIZpbnd9RVn5CA
LSLWH2XBxqHKrO7pI23ocp7e/HSI06baMqrXciJNMW0u/AcZFbNvxde0g+vgs+7mshgSmXZSTqIr
hr7amwOErfW/0zdnXgGxxDaoqYj7We3+/a/d7rtZHQ/e/kswEW1+TPGOTDIzi1rBJvIaYIRor6vx
O/Jt8ANuS+eOhx0il9eX2/gsEySZ9MlDODePgUNR/QViJ+E6z/ZEGHtu6V1jta2uYGAwAQ2gKNgS
sL7TSw+WDYfsTS4NhIBSixKB2P9oB0Q4yW6HZwHcLVMmE4inxjc88x/J9XKH3gDvs2+Bti+xIvrP
+Zu+xRkX9SeT0apxkkwMCsmCvYgBA4SSa+Fw+yDhzpvZPRUnZKWI8cadviN80Mr9sTth9kfK+OJy
za+eMYBaaqdpW3kwRXUD6mLplRIGYANixVs7f5LE4dNN/UpaUH+tOp43fyqY7Znkex7rZI9Ou9F0
Uevcot371vb4jmKTbk3oxJ7XRyW5BbUj6rd3JeFuK6FbAyF/TKUL/qCW7RdN+nfN6rFq6NKaNE5o
unTN+D6t1rlm1knjr6BmY2hgcvcdS1z8obYJqjWvcOXoQTt8AiG3E1Rt6rO1zucYAPnn9QXkOFIq
PbnXCGjFVpe7zAJEbWUfV3TrYctsaFjX2ouDRDzkSfFJQZx+pDh/T4mz4zFU65Z91aYvQxvl+kJe
8n5P+Yus2NuwDac4lXV9YfjdYLRUC3B5lL0XOIlqYdxZHu5D9mwX6QirbgvZTm7G6axoBzvD/TJd
w/n4+1/rO4eNwHaGju+1jDpuBObyt6SSNbooIH1k2qi5u8RMsaEHq1gCgAfba79I1lbONHK+uDll
9h+cDi6/5y9O7ZNkvg/jnPJXEYLLzA5WVvtIwozxkHQXcmjbsg8M29MBzNJM5p/6HvalE7UbZ0Cn
gFO8ilzYfvYQ8PgULT7ppKAsS/5CysK2R6miFR3mwJNuX61KUiMsTkiQzm7fp2gI9JNokzNa1Gak
rYi8Eg6p2BzFdJUDogAmWeltaG8BJCytan95DdbyNdAMnrj0FCYAmjO9hNemcKfGddurA1Ybiltr
DOy3q1d9Ffntay0ZH3f+mfkp0L0GDUtrRlOMyQa+reMqmemmeCbzU1vZKPUgJKRQfMVGK8pW5vLP
3h9eqQD5yn6DzcGYJLOOVTHyLKHaACkoPjBVOpS9WGd578AnBoqsPb9SbrFVSeFqdRD/pbPHyGHa
sYo9ueEO/esqk/otDNGHpLHyME3yeV36fD+xtF0kZG2ceenRE7yDHCciLioMdiWkfEt9/v/b/X46
J04X1CLnaZ300sQrmk6RA9dP1dYpztPtX9WpXhudPoNd5uRBPBpmC7fnYrGEcg1gRrtZyxRLAF2q
GnLGxq+0vMGu57fVVIlKd/pRUO+ogjOZpoGhZdWevefOPuHmSdV84M6P5Eg7UYVJf37nwhOaVRcg
WdRAWqfo2iS8mHQe+CFRngovk2Xo2lTpH9qobAkPoiggPRzMboW+eeWrGuGvuqVaDano+mljBtrx
LDHUBJsHrmfIkS26zncj8Xxy8AZ6gFh3YT3Wgx79ZiL/BtbepVN9hUXfKFo0jyTSil7xMZVTW5l7
Lhs0qOv6Z1UPu39hDhhwxKlpTXryS6v4qTgN3hQv6t/c2+XJn+Qqk2IUFVwSGKalZUm7R+nZe0MO
BeCTqVX7kFaAa4M9voBbJod0Ok3PZel6N/esRKB2btRiKlTC1PcEqJfqFeEOSscxF69RmEr7wwMu
bokFuou7IE31VRklmMGRtnSaRiN1unXUS//hvplJx5EOwXHaIsrknXY1WZkg5T5B2Up31DgEZYqZ
McR0Ke43qbnCUV3q0DjGXO9EBsHFhW+f3PTd9D0u+9g8RGYQuiCuVp27HRtx0RxO/oxj+Be2Dt9o
kRs41/N98rT6t5eHge/R+NdMBMDhgjbN4mwLIVitnXk1zzSeOID9EuIZcGhaXZFZ++9Q4HRqKo0w
0TNk3kdZbHmMLGcKsEGiLvmfVO5+92DBTCoh9aIqKK3z+oEWyiJVdseVN3CDnCC0IMyHAtxUvANB
DC2pxdw4oixI1Qa1fuRo0R5jMSuayZ7WRV6tEvk7hHvIi+GhWZw5g7goAjY3BNkU4bwL3oUUD4ws
UUYFiiYLGzEEmS2t+nf5XW0Poex5kuMBifHqPe9cqSECRuLv+yuoZ1uMM0dizNrWQ6F0Sl2o2Xp+
/EuSP734vwYvE78FdEx+mr3mEillug/NwpcHQt4zRG9Oj/tpfBPE0QIuLL7GzpjEY4nB//zSTysn
iApNmYR51NiXpgPGPk1ijgltrkGvflOE/J59QsloI+PR1ZVhBucR4NbjzS//m/z5WlhDGVDTitI8
Venh83zXat7yWBR9wiHkX2ZDuSesqhYAtwRjnfqSj+mJaCrRdYCa9kUIry4IsKZcxKxk49C/BgFM
1NoRykEUHqsv1tVRh/Nygqug3YKcB/txlxPi+VeYqs7fXJXDtUlE+OWKv8b56BhTirYOtWdwJ8K4
ne1vYc08s8Ti5h8KAQtxDf7wR6X9AHqlgMMrBe9PE9q1OO+ZTgZioZ6eJ9QNBFZ0DaaYtT3be3jn
ZX6m73ipCHHaY9IHign0v1QdX4AycZv4sXX5rMYacOwkisxH2vQDza7m4HILWjQlbKQ2+/n5vCK3
HqyQLHp+Mo6TLUQNcKh9nsF27A3Fx2rkzYEulC6eeTpjYoSKVwEKrINaG0rwhGnnmTlnkWWRaB+P
nmjP8mK7GMgOguC4iduZ04AT19zFPhdOeV1T0ELHoUXSU0///lztaek9gRQ2Qq+aUszvlzwBNhl/
RKqKv9A+hVKzXjzGfIamH/YCGPYhfgi13GadNQfXk4kQ8vgRovCXZic6fHDa447Pl3KAjyNoC4BJ
EyMRsl12EJwLE6x9s5k5N0PS0xKIoySe86/p6uHSTT2otxpZX2cS74YTD6pm4kDOK4PEKvem5z4l
6Su9JZZ2NIrD9fgD6afUnr2ZjXZyJBtCfpZ+i4gIzsXEfg2r3wacrFmhMu9USAoWUQ8EYDHdPpC0
scYG8F1ZEN4430YPBMiE6XKN4LbrDAbgLQ066bFcuXssyUkshMTfrcP4swb2wiDabyWEtc4yeRE3
6iaSllRYRFwHKm0UBCvhX1/kQznTdGS9+Ut2p5Fzb98Fi8Lkhg9b2vabJo8Qd0Yy/pu63yeJ0syc
WiX6RTpMgsOkV51egWp22SbKtW6p1Y2rKQ6w6Fv43VOj96yA1mTCmfn4XS/b397MFMtrDanBYQTK
XmkVDGcnoUrH6fzXwMmw+TMGrW4O42U7HvX+bg9S/2HnJWCdCCED1ohKf+gomzB8ZESDubdgo9nm
ngHetuxo7P5y73DDLTiqMV68W7Hka3aZNHQ3zuXvCq8q//f3zdm0HwfutgCgpqH3d7MUO1prox0a
dQVibPWNF/VQZ/RrjDugLVYPodBsPADGhnDiDwrYizvynUVzpR/zLsEN0xWWSAOfKRgf98mglt2N
du70I2IUton11i8rfDTfZKPBJxaK2FpK4y8ku4sYXBygRu25FGUWQQSAzrc7KRiA2/uYmXX2ADkk
WIFYezQyEMx/UqCgpT/rS89PG963+9l8q08au5xo5AU6V3BrDjH0jeO+KuEUxUyM4xVx4i/x0kQw
jwaJlOExGDQvB6/2M2RubmmOYptH1ZmNLfUFJA0oq683XzkFmyE2naMAtx5qFdH2jdCB1FLduDPv
y68dSmsqrVh2sOfp6mgTPnwdL4a/lJuG1qxarPNXiaosR2+gr3MaSjSiCJvlLrAKQgqI5Zch8t57
ZTnQzffloac1CTN+QbOO6pl5SDP/GuDTWBuOyBaM2rLmvaYYFEC2JVT7O36WYaMTLq7bTJnBhIgV
TIKs7n5+mK9IJzjrHIoBHJUDct6gJFgGC2wAgQw9sNhFCQTVtaogl7FwowJXZAlWM25JwAEUzpHc
cz9iQRPbPq03Rrha1qsZn4nUKMZ8CgPer/eAuBMDlbamCZYqXva5j0rREe4uCska0Y6os/7qoJO8
w02ZfCgkv4NfrMGa9Zx1CPs4gzYZGPtwXjdRtFD2mWc2aup4BsMeq64bXXXcj4UdmXPZlZx9GvtQ
XGEGOt2hsvgReSzSRJQIIxqAmXn4oXZMowqzkxB1f5g6ikIRwakgheGGJcywCEtTJSGdWT7WcfcT
4a7fkaPgRxnSwtJvQV5ewRFJxk2Bt1BV3h3Coj2BhVuvhCIAtb3sfH0QPSajKfCCOwnro+VbrUVz
9wqN3I545js145btol7OG/LvPXW9dQZ1k9zi1rHhBezsn+oxdPPu/VlrDikNzQvyY1Py6BSxKei1
9r9trAhjmx9Winbh7+XSJxcxl3t2HaB4S7RgU0Neod9Ji/IqS7cbU0kLATycW6IB7j8q3W5eIcvM
7BQrJO+nC6hv/mUQp+X94vLrP6zPOWYP578p9fRqJV5mywgbEF51045/jFLgYk1oNwy386Du1ywb
sDwOdz96i8M7lSmxqp+omuB7jU4omi75kio0bz1tR5gnmV2Bw8za0s6rzG6sHfhjxOZXWzm46W5C
ofFjE1CJAb5gABzfFcg6RLLLU2kriaLvxAwV9GgXRHm40gUjR0bk00RkRluQIpf/4LF72WYGktrL
PuPY+pkrYcxbOYbDdmVVN3M8+LYxzr6tFLUjoF7GQUKR2FCxWhnr//VrNwysX24+PB4pl/qzG2Db
ylOAn0yxNuepik2b38mwpNtAyCKG5hu+6aW2uLQ5TklxOuGhGJH9pE5uOyHwFmQDtbGQrART8oHs
sbAREDec1Xo5EpgbKK8VSYnpaXmnFaBcP5lQzTvaRnwoiyqUTFkxfchGICi6CWLuYvIIwEvq17Q1
K8GeC2MnxTAxYnnngrC1Qa82gEJDt8gZyDzqV9pB+CgGnADx4Z0ETwbGzdtgAhGOQcP0fhz5zl2L
AInMPFZl1oGmqj8kToHUwH1L35cxmL9Uk+LEZ4EngpchAl0tYilnbpEe16BR3OGrk2JcAPBm8tWF
ozSA6Qt2AOeSy4CExJsvqUgbP84PqsXP4VbDG5c9BmBBwo5N6JTxzsjGbJC27mQRC7RBdsZqxyQU
y5gBBCy4ealaooio3u0PKtuazT5SAiGX275n9GgEFVYDlspWrxCALM0vY7IFjAVIe1BHPdqZ5/3W
htyUQ2jap7RMRTLqj/zp9hyiDraqlaLvdWAax08jAdP9hzdXnzZtsYK7lAtrGwrCmUllPUzlV9Ah
//jC9rY5I3JZ60CjtmSB63ZBHe47etFU+SHPOhh5rB7G09wXGy/sAPKPglgp6sdNKmwy7jgLuceS
lC+AO00NfvfuFHIPVetZZoR7z4OH5b/0GQ4IPjDPpYyqAaj9ChbJmOQbFY3juilHU4s6ECkG2HbY
9RbGGaFt9WNiwWyM8x0whZlRtOnR4wQ6L0rSq3a5h9QhxbaOwXyF2Lvvx5tfVVzLdV0RYsLBbObI
SuAvPusdhKuEsWbmYEiprgtw/LMHV2nzCnaSP3ul0rdntc5CcX9cv8jiLEEkZIzQgbD1lI8BnaIB
hDGr1FV0zaOWW+DVfaELxvxPzk+6GqzFky6+RRo7nWhBzVZEP+4utIl89diQU/SlpZI9YxQxlOlv
pZmL4cx6pDK/w70yd5ouGvAKXjctLVFboVCwfyxF7rIwYrdMBjVCvQ64en68NQMi9BlH0acf2ZqJ
ZjE2h22d8sjYuHCfWVk3M9jxf4BUB/itBisXHjE5sqDT/Meng/V7Li4shPrTWuhTmISgnZgMm3FJ
GeWZJTrI9/fBdGjzCVhRoRwcJUyS5eikQ3Ss0VLJnlCMUmP8JTkt1zJnJiC5KTnpc7tw8Wvp5+Ic
aSppQr9T3SnzuTkNbk5FSD6pArFOauL2xGfaI+09FQdWz+/ioPOj6OnAkbf+Wie4sNJEEnen56bc
D6JCiFAzocLVuuxV4ucDtCxNhD879zmqx6wkPbpGQcQtC1UeNukpkrQj+Z8Itex8N6iiMWb6/Rrs
joNKGXa1TsOVZnK+KxsNLdPbe2ENzNPXzrUQ0RDtakc2aUKE9LJdSeZEiqRSd1ykvgTzIIC/5toB
1ByVpIhIBUUtNkMej4uPW0hrwo1Br5fI6vp4ol+EAu3zAvYUn3RgEMT8mnc/9L/noAKHZhKfEsyi
TpArq/KLCSWTp5mlXUcmebvCPl+kIy6+UJniZo243DRsWOOUDtaJmF9CS5cijvDGd6PkddUqAOcj
RbuLAW02pjA2Uzl9LtOdvtj+mPzq4amWVDoRFbjqdClDitz/8qcMRQnoy3KfRU4u3PlJGh37GT1T
JBdYKzjD57PFRrK2vpqtHsRJ24PYfbu7exjSLsav7MLSlVMBQCGh+NAOaN+BGsBCDrMonEgE+6F/
CTmgvVgfFVIdRuoDP62OnaKq/0o0zIFIxarm8PyNOs5BOqyCbneYS+2ku4bsjE6KWBJ4gBNUdH2d
5uJXtoHkaFBRYDkWPDWYrMvLR5QwVZjmdAxfiWdsICMlXB+CS0viONHDRpbEg7WMeL+WxRgGlAon
D/0Asaf+kz3SmZx5OWOaseZDLBcvNNiQvzFWjPW73JQbhTtIZS7Krc/4t/BDioNT/yZYtn4WBiQw
VxW8FZTBTuPZCnwG+yMY1zVKl7xezFSAtiYtDOVENgnWsrlkFBtsj3v8O/C7t8A7gQT7fe827grC
+pTlkbUS9FmRBO1SMwijbbFpYGFmO6+Tfbs4P8PtMU5gHzZ5kDA1+S5ah5dSd4ChwRFku/olsxIo
Y6y3iE3aM2TdLUS3cyc4E2zvMIu1FE+7p7eBlVDOCFlGHwMiljbfGbbqGdjk8ZOqq9vaBsEc+pjj
tpGktXwdqvgq4PFI9wYs5QU6t1dnJo0RiMUN8kdbciVNNjTp7LgN3w6rnfsWtC5FuAf19CzU2X1g
A3hubd+JEvnfjmZRFT9XE/kVl7R0rn/sWxZbHZ90h8xRXJEzrmtK/hfkmbnffz/ov41E/SxPze0Z
DoZGAWE7+DOXckOtzXzKhOQvMIO5w10UnkUChV7ZkHX2E05b57jXichouZflTEPaTdSGbdACdXju
K2nfWl3YIEi2OlK+YMd8vJqWAsrvhiAfnkTxqZvWZ6uTSyKz+TVdYERXf0mwctpFkd7XSGqUAQQB
6wZUYLWadETT7ujv1dZjufZ94JnLfa32W4tCUj2ASZWdbxHB/fAMBCWruvMfWJ3E4lR079C1z7JC
G67+Hh1SWMLSWtviET4hdw4Y2DE2yLF1mx6VILQtCoX1ZYXNIo0IlszaoChhPPEIYEQbXPg7RBPt
dRSw9Vra9PWikxTaRaP/7fxwsS+pNe4mnTXBg5V/OqButlevqPc+k1PINnlPVY+XY5+4yJOFwQsm
cJ6T3/TYzquiLaviJkNxO7A6TKZSrgalAPxlaJus/5x0zkmgIayROa63Kc30s2n/or2+rmmul7A0
C6UaxWIfOR2KCPJN1Xy/qabBnaR4zhYUemr7PZ99SXUqhU2+t61K2avgOZ8unF+52knAbu+uajKB
oyyascGL0tZ4I2I1T5VtzAm0awqImzUrz6Mdl8roI+/CG5t5+EFaV/OrTHyKxIqhmgo90dMDSwQe
SlJwe6nlv2NXuI13P8GGNpAZJoE46agaIKyt7y9WRXoCiuZubB40j+21SGj9eobU8xDqjTKd9iy1
jvTuSHItCRbxfEz2+eQhcM9bziGAga/fhbW6S6wCnJHFlY074rR6VR/sjIUpqVFjm533aUsjOM2J
zsB7+5sfSOyTtkD9XMsa6WSHG9nGGe0yXDKyr4iVMUTJuEGwY5JS3EVwGGhl7L3nuEjxSn1veniP
egXYAEkhKnZRiw/MwfKRh1YcClJ9zL3q/waHwk3b4yyrNn9efBEXwfumJepYfRb4PRZOYqWXAcd+
vlnLrdup2RswimHfJ1n5GpCudI4Lm0HsG2ZsAcH5s//ikcInWjgpz/7zNP11V3zjHOPVglWLWH1+
HG6I2a+w3aqe7seR5JlTSxc7ZDi4I81RQQ5F/i8+w1TRKLNjD2oWRhP+U48JlWQ5LDDfpMPTKHyk
0DAJ8iysGAmyDEhh0DIMXdkcGSkeIDDeUgngRRh4Lg/ldiJmaSu4vRupSBC5XxvFahrfSDCq68dN
1jKkd5iprSLy/JPgN+RJPZNYsS1xMIU4VwpMSKmwphe8y8xVRSNoySXHsCPNuX5grf/o8t1P+HyZ
KLCcArGe1ABntsOujD0qNHhb2LU7ywTvP7YJmQDIznnXcpWWJiyftFJXwZETSrAF4X7tP66ARV1P
7NlhM6rPh3yg9EtYyTg66A9ihMUNT+Gw15F3vQKYFNlu9WT8c2eIpwFy3aHRD//EsP0PQoDxmIzO
A9LLG0VEaI0kZrmQH83pY82ea/aQGu8vhMrX4JtJPlKeZ/QXT5QEEepNgrrQ8WcwIdFit0SLKjrV
GBlto7/U7dHKlIgVZOVB1380HqKXgq6ELYzz6Z8Br8+xLWekNTmM/A6fyv8L5vSr3JIExeBVX6AD
2TcN9pPG3fhUStB6MCFSoptTuadQU849UOaAsqrxW5Kqihk5FHq4HpXMShKnm7e132P1bmpWwU/E
V7TDUYlY2KOAGsLpkVOkfuzxqBeuY5OIjoQ9PD/7cIQx3CvSn3zQsIHq/5IJTrC0+tKRLzE3De0M
e8b3D7FxV6xibm95lrxnNhzEwaAhJScY8T3OFs4SeSG0bERrOOmaam3tigLO/KpJW1SVwB9Q15Gf
AieEXE2CCFAGkhLK8TQsxtxfwpz9nLB9mtpEH8oHtsg2otlcdWPYW2YKKEqCWZqsRZ12jI26rUa7
vxtCiMMsXHoVSz3kNeP0ykZ5KmCld75KvQXz8VIzAwGT2Kg6ig0em4ckEFbESDQtrb9KJz+E9KZq
pJUR7ua7L+9a0Fs0sruFxcMXpUqbDUkUJ0vlgb/c1FYmHXeFpKh3/S3POO+JjVNTAOPA0eoAYdTj
EKSGHKOsfO2b+XGBb/7iNhKn4NRxncWsnDsSvx7oSXSGIuCHG+/DrGObngVxpxx6hljeNmCli5ap
48F4jeq/AlmEmS3GfJUAMfsiNg8oynzmCfyU+iHgrSIP2A3usypHJNCbxGu91KJLZMY2hj4d3ap0
GbXVlIDII9KXWvtLDeVIN7ki3W+Psrii2vIQq5xeb7J8CPBQvL00TTU+5RryiwoNDsRveBdnVNwy
B4ERoM14NGlx1eyTlDh3VYPRO9O7S5tUg2oC/0b5EE0/ff0phfXg9yAJCjpGIMQn+7DTwOkJjtnF
XL4rlIfObB9WSSeV5JCjhGWMRplbeQB7ql8RmU69v++ZxL8/GrKqwVoOMEqiYA9g4sjkP9QpK9Od
x33SfD0IW47a3tZcoE82j7ijOs5jFHjdjnN8WxK0iZbJPYxa/diKUpqQkYMh/AP6AEb/LunFiMdF
07ronRzzpd08ae0pW7sIQamckoL27VlBhfFmZE4v1fXfwKsXGmFOkLfGkcDvqZWUOCwj2VFCaLfI
StJWN4ZXSJobwXnXap6sCUyQ8t+yJs/QBBCvjA7OkP1nI5zKSWsewv1DnqHybF9Usmvlb+Km1q0K
bxxXrRdmYdS5KuLz+9Mk+7DZIxPshMcX9EXTfOl/GR8RBesvGGcTMKg0xHyywLp/lqkFkJ0pEL+R
yHz9bT7PnQVcm5La/afgoxLUKrlyXH9ntmAY/ldsSlPGZphzsUoAi7/eYau4GsZKU0Wy6lpf+rsb
aV/G004QLVfrdLCxq79Edw4WgugrL2LDfo8X3wbM/N8Kh/Lcp4j2+o+Z1carSVhfLEs+1O0PLg4v
K/UqJB/0nqBge0U/7EVTIOtpF4nRRJwWlqHkp4WnYQ3EBcKVlZxAygNxp7RxZJisovgTuF4HAxQM
enMgjnjvRXMUMStSDX1FfOhbc2riijkKPQinnFQf2HxVayJ1O6kdrCYSpXO9ekP9podPWOd6a/sO
ZsbivwRFNPM4hBHcBf82FNZzqKdDSCj0DDGFP+75eSzgIcwnznuObxCRapHXnTVOx7xJLwI+H2B5
FDuPgNy8j8PL2iaPLYFNYJqORX7Aw1kzIpW1UkDIJm5zFtn6Ga7Qyo8HZhlgZdPjeSb1PwhxcHJR
t5T8qxZtzptZkqydcJbmN6T4Tms1CnCnxGEsGjMjOTe5x2oAg1kpqC8va4CmNXeOrGFxBnnQWnP6
+t1HFEDihpQMrBzukuvQ2qT5F8eBlbZq+kPhyz+LW3ruW8eLB7XaXl0zwRTLaDi2IDRy5Z5QUlxZ
binijH4CXhHokIum65aPEu4uP+vhXyJ7N2FhP+FVJMXs4l5xQdBx8mJpE4oY1wQk0yJ2bJidBObw
K/Q+TBEixN7uOTHiAwLNXM0uVO151ixcHb+XwCMpZzuR3+flegd+fG0dewu6nzJjlDXZHl2Cl3Wq
bNIpKCar2XRDLG5zzyRgQUGuUTD3C+TIxmD6ZrOPR7ctlbj8HMAYeJJekSf1S8qL87aPT0foXi8R
o8SxYoNFD9ziR2uitGamyxSo0OY23UVgoZKm9daFTO13sNhqnGgUowqi4dEiAqhj11BsxBf82Ro5
7VWCJB1fuPCd9whzXbLGYbSeaoSJw+wptXlVjlkk8Lh2ZPieGioeCjMLdDALb3NRSlUxuQrFkUFs
VHaMsze1uKN3YdkIKuGqX1xtumMDZj778EQ753iudU4GkuqnSa2U6+VsmpUaIPVBTsFES4pvpyYJ
ZBl2nN5GJixUfcr33xttSlIkEl5mBDNry2Yo2QY/r/LMfU+5uWv1vxSA9LTzfpciUJmOhioI8QZN
Fu+kF20+n/F5Ad4UNCsnL7jJetD6/zfb/a+xPSH6udhTAZbZyLKhLhqlirrSw6AP5rUUza2sG30D
EHRIKoVaKdpJGHgF9OdZM44TrJCcp3VTSpIwJB4c5tLjTGZBkbLP1nlzHsveSP7Valdpax7yY4nn
k5ERagvnIdTRh6/X3MsXA+/0fFQP5ykG1rAVj5cIIe84y4eprblLqjJQtoABd0oy0JiODZLYPS3T
961sMYzMHFrIWnLgeNJB7AI+j8Qtw5UJtnLsUT5rrkipcJytKJxN4cfSQBduOV+B/LrDI02Xi/kr
3xgDYWtzi5lAJZv1HTNlaW2BAuVNf9Rnbufvh4WHzouLKVaVROtUlwG0E3jBzYQpFY6TrsDPNbKO
pT7VlB81PvZa9T8pgbtRZoW3dScVkV0HdVdE8R5749T22kDEYdSJVgXgRpKSqPHmMOqqWooJYLQb
56DSMOYoQ1v/XRTCGS5hT5haCM053tOMKy5VzjzV/ksdCV/SFTtJbuowvARgFJRkI85OVKwG+T89
67gh+FfwoalKNlsaarRzvtj7O0/lzX/3ioU4itwsUZQhbynjpFi+9rKUZuVdp+I0AqLKHtxAfoIP
qZeZG/BYPpbADHRu01/EJ4gkqneAdDrS8p2AGko4sxkdZmFGORid55H2pPqxtF4Uo4JekAhtH81X
gVueeVdCvi2M+FQSV/Rh69lpO5AQpBZoyc4qtdget+Io4FLLPLR+ZfQSfa+DxBHr3jbm09F35ILS
e0SC1PbIJtGAARBHmOjzqjupuWMyG5FHHAN8wc7gdy86++5r/tEVTe8l7kZl/P27ynyepfBZpN+w
EhmVn6bPGMZlDkFtjjXamvu4WNZzJoGx7aqO+Y4kJnEdOt5k3uPTBrz6EsSyRT/okpDYKRpQQnqS
G3c89YcXx3VUmcXiaPIxTztRLYGql5UnRH1WR09sFbiPUAP07RBgZU87ajtDBeHTp00rxOzheier
xjLh2GHXPX5WfWw8WXIMjJ8ZO0+IXD7kycYm9eHh5NgIb5Y6JoI8HajFd/pv6bww6N6RdtIW9fqT
4WOhcT/1R7MiIzTNXOuDoYlbhyDCO2/QSn3g9AD0tl67MPavQVroKSVr81XuceCAxCIygn1kJROW
C6z5NHAO7k2pCq8T1JiUhcN1Aexbwhz46S2+2LyPz6vBCaWvs6O8K7tFYdlbA6a+y6/cbZExSnN3
G9Fx+k1k1vGvyrfxkCZ711oGpu3KHOVkL2nnOWqIpdhnxrb8KVJqIVVVjoj9YUlB5QWUWjyigP5Z
IImBQizRArkSG6sUaf6GcAigbTIX3Ut3W5sa4a8e2ZB2kAsI+SYwm0a7Z5mZwPJfrzf89kSLCVeA
EPi1k8BhbMgxwanHea440X0usOhBcQRi3U6YetvRLnJrfnY7PkQ+9YyBe/g8PkNRnw+rVMT/9kxz
b8FNuLZ+hgNbgdI85dRn4CvMgfAh0fuC7pzNiS+/hDNqLgV2QZPUPDxkBCNkhrbcV1WZT8Oe6Dp+
BMzh9nXyvGJlp8Os43LROms5LIdUdFfSifk1hpFNvssI2uTEZ414eOG1yboA1cdpK5LiyYTx0XgG
PDtySsKQVXP6a9pa4GBI7uDOoIMiyx3RofJysXiNb2PWAKsv1FZOBqoq4IqIsfSgutB7ccBs6aLQ
hnvx+Vc6UHT+YhT6MsRUeZwreHlqloQ3oLmG7XfsgnVZspDbmChJOKPU5mLlV7YX5CMYEDO9aAN3
VOT2iuBqxa5aSGrvZOfADam/xQxcf/mktu9t3PDelGAwn5SGMb5VdaX27NNVQ1jDXoo6W54YkkfS
OhGyqHSZIaa4vuKrvzLb7A9fV3naRao/BmSyguTmGxgpIvV91dUs9R+PMOiMcwrkUx2oCUTSEhqg
1rgnVTFQYMhAQfEtX6jXozO8F3mNNh6fm8r6F7Vyf0odB8eEliYBy4msQ9SwOqu7eXEVJraMd629
PB+xZ82BBgV0dF+cmEhcOoTtYe570aRzTVgBiWsTR8qVbOaQJLK6XA2pbZZa+r/LuLRYVqhX7lBs
uBGfkHoqoqH9aB293U2kuJOVcuLGJNI5Ih7YuLwvqCC/4iJtUz4RRXuSuUDcvbl23fTrjaeYTQpl
x4HULC7v7qVDFGjOV7TTIIWy2aVP/uewzAky3IwkUd7q9AZVQpRVsK2upEUFiJ8Nry8QdMjwqv+e
pxfw0wfwD8GROLzwzPZFCOnZ4I3U0CPIO6THdoiveYvoTupdz1/nbMexjk3sOSvmF7dcbZz/ACEW
9OlFdpd8i7tulDthMys11d6n6rRk7CqcvaNFBOlrrxhLb2qG28CZ0ljKn9qPAHZy1dcUkUT/xSMM
zO3RAX062rhyDAN6LrV0hTxoHIw1yYUC2mlYzPVf5uzbjuciR02WDyAefA11Le6Xp0ug8TRz7Rx1
kPfXjr83CtR8EoYEIEGT7qWSJY+satvro7VNMKWmCCio89nQwlcAw/k8Uqt8eMiZJFV2K7OzoQn9
/cphO5JF6Kf/i86dFxP+se8L+UuhL/0pwkJJHF+H9GGsYUQ+AgBixZXT8T62ULgShYm2TKSsBHYp
bZfDr9GeINGxfLXRA8+1ztM63I7XdNaz7MOhESZ+AK3U7z5AaYiGdRIPisWz7a2HYl8l+ATgO+sG
561Rc0o71B2Z498eGT4djmSNYCP9WUMnx4Ndbp+R4qjST/4+/kCJai4CGsdEbsp4zOWc9cFe82H2
GhLPsOAztN/y5IqtRcur7IKgNJDCHFNca9i9oJzePIGlh+9eChN9pctBsGtr22IDwjHFtV52InmB
1ZGr29qW4ClppRVSSJhwtVDswrtMsyrm83g7bt/NDYT6LLJjPHGLKB3ipND6VfwGNnELxew4IzZ3
1Nm9I6z41bzP/7mEAwoZMp2SiS5q/B4DSRb7OdGNP9cvBMD0r40pojvdjOpu2iTutLljm7+PH83H
Cgleel8rLsau2GuNGs3xtwXafU86UWxkhjcp2Ur3AmsXZ30EcFiqjLDEJHCuEqhpdu10+Pna291c
lJ/6LWdFmVrEGwd6UYGTKNE9OhOTyiLMYjBaIPrEO5yRsopEGBtiH3uf6xAqLMHLfce2GSk/AUjh
sioI98scRr3+so/0bgVkIEWYg5jv+KqKvl1pHaG2aVXUxzagwsBbZg9GVsoVvoqn7HvG94Ywmd2P
mYF6LnXpiuKKTtTVxm0IzCJSVsv/rgodOVoVrOICz/C/eE7S7ljwaTKsFX28SIA7CjBYjzpZ5k4m
movuLSQm8c4jYm0rvrqRNXmxlRxd4qUIUl++Tn4SnuIPSAmRq+8tTlPN80rRVDOeSUgV0fT5ayrs
mLD3ZnfvfhBbRfAHt3/GmmwpG9LIy2/j1pA9ISwlDQjOwdreUaMLbrwL2AyfGut20/MvISfL8b6E
49zbIOYivWhYv0NVTl4t6FKbLjRZfr4JFLAkn4Xr3W+ACLikTZbRue+GS6NwU1kiRYTcgV7fMm9Z
PorNyi64Ka0+M0eKG/FEoofLvf1mN59td1jd72ek1/yT55qahUnrRssZBtjeRj3Jhxa/J/Um48X6
ofRj6r7osOzv6DrhdyVOoDTGllIqyARhuPfoV9i3DrtKvKe2E9hceDD3QemrwXd130O6yZn5w4sF
k8+Uu7ZXIiRZ7tyo/e9qmBHlnkcc08Z2vRX+5B0hczhqMyh+rNlaFUnJc3sjGrUqZ3xNorXm+BsD
RlsUs4O98P3MHevaqK1/ZczU3HUsrlzz/WGwvMVC0eB4c5c+NzYKryOd26FUqmn7LqU38A54AJ7D
vpx8cXRtcMkYvHxaqeiXa2HQW1sxPmj2l0f/JT1Yg3w5B322ScLBwz3t/4eBjtzmVVaO0p52BbKb
RoRhm8Jwwkzp5o4wGzQXYhYpAJeYuIyk9E1P2hO2XBzwrSp/2gY2F+OHzr0defdNUrnN4ttpGhbw
m1G4HoLA0mXYhYWlekIfbFKcfsoIvu4c1vcapW62l/SEc+eqE8p+D8/v9XP4qeryKbhjIAENhdlk
L47sFG/d5UqbqHm2E9ZoxKDbhnkJJzNmqARK5qArNvelnu6Sss9ni0AEspPIQ4Lz5c6qWG+YKE4b
2o3Z9/AeJg24KlNUjLuPRRU7qDmD0DCWsFqB2XMen0tlHa5p8tJ2BgqKUTo2J4gQp8qgkv50Lvbc
QejKUx6dSIMI3dkJ3ls0tu9nidWozaT2k3lgZ3d++XzZlWvsgW1uXyr8TXGVqIr28Pvpp12emLSs
3UVXk0QVvPp3xEbwO9hsjiI0OhOcYaU7ZRmSufe3fs0umkquMNiE4GrWKcBF7dwh13yMhZytN5D4
MixeI3b/apCEEU8eVPWbsqyaqy8wg/HPS73Bugj+z/oqOFwU6YYK1MZTu2eqP6ZpyKK8FQUakt4g
TxHjXg6uMN4XmHiJd6hn1G337bp6PUSVoSt7ozvLMq5woq9NjI5oKL1TgMxUYbSkHVRkpJ/8f/wm
d72RrZ+8AqwpoEMrEHplP6mwXxBg3D1asMPlMZ3nnbc1A6H2UIG22NIbGTj4aY0I5nqdD7Co4MkC
IjWYTet8CpGwzuyJpWjIR2Nh6XTQ56pz2OG9En4i9UAwNvl8g8aVQmxH8bzRZBKNb0SzwaPQUUod
i1yyUsF4VtFuHn/MJrf5AuH5N8qeZIg5KBeKd8cxcdDkJbMJlQGW6R88Ec1/QKUiBnECEhOgKGPX
aRl48sfLbG1numS+x6Q1mzEZ7wc/JKjBc4jntHFdd9Vzg1SSd12hmKJ7zurN9BKxA9xzzVgXNbEe
+g0geLDGU8w+dvChCap/NkwU3+ndxe11T05sPb8Nk6DlNhFKruo9tqkHn32hEM0iGobIDyCu8zpp
euSGySM+XkpKEKUoF2++fadHiZn2jSoQDGQGbsm9oGiZ0OwvAuFzxTWUjEeUXJs9fgQwHUemCQiF
23hQEQwDIVgUARmnP4+7Ju2rS9mOwM6vKm+jc1/qoqm4lWzJPo0whX5zg5OeJUp4OwFYvjespEcC
9xDp+Ts2kCLgbHRXMTa2l4nGXOgLaBX0yd+AHwVpig783YaWpHVISiAZ665z99w/bcIUjsVJvC0F
6VNzPgx0UPcGzfQjcYVlcGX6b7fbaM5998rL8wvXPAC+7Lq9iinUEmFZZI/SlJ5fW85RR7b3TgOO
+DW5dzHPlqkPIAEXfBqt7LfMucmbwmOI2KzVK7S1ltUO27YvVb9aOoVkKGy/SSVF+MpMeY+Zn8RP
+6ZUra4XD9t7XihqMTKX2IYkq9KC3ouq15S6RMNUlfw/NRbX6K6ysjjNSFyYf/W6PJL8TVD6M3kJ
CkurGYZpYWT7LYbKd7Ir0CDcxJNyUmK4xtgapJYEzvELt91wwMhHSnup8arJJIfLHHfElW0BxkOU
XRremr5cCFqDeUTC1r6YsQnQZ1gSG0a8rzaJfMI0CtnhzE9Bzah8rOtO4XnKZxcDM1WY5sJCcmT+
3opNn/Q98jri8xpza1S1CazhPlfL9BBrFoxF2/ziP8NVpIAQyyrOEGx75z+SJCfuJffHzmnkz9bt
nOca7mgHCT8UqW/lXez3X/3ouaU/ycPhcxgF9PEnfTMRkwiEJaK+iA10c7HImIIc8siPCTvg88ZG
Lq3N1CNoUlkLgJ2Yk/0t9h8PjubsE/d9Heq4xF7rhR/7/ccJqcMnwmXrYlf6vnobo2OrpwyXJzfu
IrjGMC9TsvotVKHSXeunN17opAqxT2za1p7f4QOeWwIOyxvJ0Y6mSlCsB57kl5ahP7gveujeNCPP
fctcQhdNNKs9oHTNJMlDQxUIihER81AA7vovJ0jz6m77YnJX5qUV9cYnP/dL2UL1Hu94Id37P5d7
/M2Hzr94ubm0qLqor7Yf2scuSluhqzWmIARmtGY+OZEcv9+jgqDioE8vVr8JacAYVgeij/+RTUyX
aG0dX0qlQn/TadGJAXvI19WwW20UAFUBsWWahtb71KrLTTdH6G0K4oJt7JAPn15LltvK3m0vbCX/
3LIgn0m4L7mKBmBCe6vuj25WdGDTeadOXFDbj5P3l7X7XuLp0OA6uaxz+Dt2gdQXbg9uEXM89Q9q
xxN6+o8wmcuZveh8szoKVfzEdJoDAek2P5CUbrQ5InEPYQvBrCpjzP8LR/QIoN3LERLflhLlw9Oy
072OP5ELWGDCGCNzQ2V+ZbDtn4dGLHqCelJ9T+JzZeJAahxru/ELJKynHaCHGj9zqd5NpOzlTAnT
pZmSIt86ap3oXKgEDAfiNazr2Sgu3rZK5USMOn7gC/znLDzdKhTurrsZ58a4glBY7bkihg834DEK
en0quExr2f0j5Nvs+HMNLR/vEyADzVLhtXjVDgkHi3AAYau2ZhXol8RkfclmrukDhAJ58Xy7sNoK
SZ0tFPCwYkm2XgPirpRtauE3BNVN8ZqhZ3Sc1pUL+eAWUiGI+ZcG0XfhjKY1NoVM+iDhP14+5VaZ
YUj3bIkvnctjnWe38zR3gvbMT2vTT0ZlUmO6o8I07FrAvrYcNQ55PWMuXG1r7UQq2ycOZemPU32e
LzbfZN4shYJHqwZSHOR9mTVLYIL5IcAkAuDgoAlrs/WNpy5Uyil9UK5MSG92jNsCPwyQPFk8Y2iL
+CJ/MwaE9GgEraGiyY1idedHM+u7LgMR3DrMAE/Rfhmtnc1x2yTiKflMOABJUm630AXG2JrJ/o7I
g06oRnhvcfd3d33zgXpwYqqng79EUW05IJewhj+0RO335Ljzasfye5B4gcR8mCBimXn7THISPRFB
x+bkJUfmt71B1A6PE1L6N19iD5hGtwlsoD3+7ivzFDM/+nfXZRfeC/zDtamAY4zpvpdHp8gqGLFZ
xqIvEHm2gBSQa/33n6mkgK7H6pvSCs0TWfVS31knKaRtFD4aG9uyKDzUl66WxC5RCVESrAv1jXoZ
K3H8oqAcxTfXOs0kESYaUozg1PpxqFlJ+oUP8bvJ+c1MsFZTWhyHlYNH4j2rQc58P/+6LKsDwg+1
KLZDPT6nZbcK+oVkAI9A1Kj5LgktSIlZ9i+V0HOYuBlMHyDYQCXIzDp7olq6trV0fPRR9SLRQV+o
vhXKSWG3Umwn90qY06N4yBNnH3uv5mRuxDeVcjv2pXaX71DfA6yi3w8IG74MjBqbfiPXqUhKNbPk
qnhX1RDxnQgmy3bnQQ6it6aZvXYGUPZcatHQRgHZYXzbVt/aJ6hSqw5T5BYk2ItUdd29xDX8K6LR
ZUP7ZVRMSfJtdPyYfMnN4ERIPWJEObs/ND18+Onn4YXj3NFcBNuffZyzhWoZ+WJUY9gsgk/Vu65T
E0DlfV2ZdPtf9G0mgQNNQkgQ4iFIa1j1k8t1TgM3qibU3kPB3Qj8QzLqGxbPNn4qidWhk8lXYpqz
LYIvyuKyBBhEUxZDOGXj+D5ts9+dYU9lvBTmfK+TvlE8Qfjhsz6IyybfVp1/1WcylOVPNb3OL0l0
7cmwYbhAHcsS/E0+onZwy5HIaHRczJPaHZqW/IdLcKbQ/rJML5QPVeJ2rErD0DMAkWMBvjg0gWr7
wkfOUVacow5YdEr2JnHCPVcHX2Q9UfG4ud97TxneMCjW/lfRFJrjiAS2cKA3f6Rd1mP6btif9IuU
3kLH/grSQSXLiyQ5LFxsryd4AwQpXFGj7FPXyDTTQ5e2EClvG3THSw71BdjiWnU09ZO1Qur4uyN7
SqnaefdUVLuZynZ1wVz1j6QL3hlf3WaUGMnW6sxL2MMhtU1cs9wXo/y7t+XnR6+AMNXrtdaDwtyn
rsumj8h5r4PRpeuJl31UVEJhB9qhtH/ZdqffzYxA3uH8LBBIUWFrW2m78WDEuLQF181njWbBgdC/
9nRj9vkB6XjhnGY681dqCIM8LVVodvUtl4DEY8v6Nf8KCZEsXD1N0qEFK4t0ie1Q457glpK8UZcG
EBmk9EOccZvo8KTzSgryNtsnh+GzvOMI1JFmaokaD2Del2n0pewrQU9k6NB5Sc2llLv28SmxEbaM
XKc9m7UlrACftkLIF+cYsDTlbHF09NpUNfNo1hTAW0Wc9iBkliLUC4l+DJ7FYsSIMsjaPVG9r3EU
ukweAI01lW0Xci+NiD1X06KZinu3NU3845R4eCuairsRyfXFDqS8X/kMjVz8ESgT+ODIlI+Uh3Ld
kriNBAT6WXGg9sM09PGY2AvxMhHWIudqM1GBXGsh87JyHBNTWqelZNCx1Te2b4J9OfRHX6fx+RAz
zfDYKKqOVTR8lrJrpDLsMCDSMJMbF8GUnf3240s/ZTDWDsnUIEDiRN//TNz+eLVZmJr2ipFEx72F
GFF+OOriOhzYpfCWI3+JczYUuQuPuaCmXuZLymdzM2kJe/FtF+kXUJAnUiZ2Q0KsxpmHOdvmc3JY
wki5VZjMYinNbMW7XB3lkBeN/Dq90AbofHJrie1OdB6aDUrjVflUM/J1BNHooz5fD6ZkpUdxqcGr
t5qJQaAaVlZwxKE+4GA3ioE84e9tRFDtdkPklEDrNTt7xkzfAKqxhJwQ6mUFhwQrZ1VnWZCgQogj
ItP8bRS3h29URSJmNu0TQoBB3bTKpKZFcvn47StxuuFVATbTIq06WF455ipJooecLzN97a3zoOem
M38mpEUv+9FfNXr5tk0mrROD0PS9IFP+D2Tt1p4EzfUqHCMYeCcc6Dd76gLO47TJcBsfdTV/eXbg
4bIeZWOkl7JEa5efvlx23DMA5KQxFRLeUbJRJ+1+DPwJEjVwPwfn8zupQLxLJHR/F2qXhZ8mwTFi
xjbcqSg6Ausr6f4UTzlhIY/xXrCtI53pJ2jnq8jsmyFjWQAM6xqBn3aZ+YpN5iGVwjnnLd1ErTvx
hXASR/XEprU7NqazK56bd+FSyC5LTA2i01lpJxVB0S5Gxyt1bflQJY/GE4xid3KFJ0A/4TALmaSv
OVSb82LEZEEeSoqPeYbgvfAaGwopsXWmHBN/WQERy/N9VnkvAUgpYHa9ej/ZLqN3S/oMFdd7HfNu
/eJwpXIVTXOI207M2ToT/S+8lymFptxLgnitG/A5fkhpJmZVv4WyPgPgpUCLHeswtrBXQRrUYA30
cWiU5+1nqbl5i14euByRVmUqcjGGkicC0g03RTrjbo0vmkzs/zBstpIjPAQDIaZ9MB6CGYqnYcho
3eJ9YrV7a9aJYZiPg52z5FguMBlfYqnr9ezLhDwqi/mRgUaKkwMoNHO4phvXQhQdmffu3jUrmrYs
NLxRFk79HQ0KKzIawFvGz+fLvMrCQhkJuI0aeMcw1u7yTxezXHO7KC46Xx2URO9Kf7sKUpKD6gR7
CHUcBzwX70woXel7tj75dvyfa562ImeSeqp5jIJ8ZQJQ4ilY0fTPTq0CDXGRk+JN+R07ZKE2ZBdS
pgy0jGtqlZh7cKQtYxzb9Mead4lPItOmMqjQfM0VWNyt4lbFwvYJtInka0Uz4UJz1scOi2HMk4fo
0QWoPHxr/a9tnQkHgaB2H0Rn1mLh8TEKIskcOSfvNqQi2R5nHClwMJESMzSKxgPtU77s1CBcB0l7
d7gCdpxKNo5O9p0/2vfL14wKZFG6MbuhrmLCOFUWEbraZWFbVPy4dVK1YeFd0+01F4dUe1f9SlRB
a+wXRuIJ3AV0Ziq+il02LK1ZZZCGlyyzrN+Fk93p6NrJuIfpPyvLVwqR2CJUjAHOoEGTXXfP20fR
R4gYWWb0tsgljwX8a0c8yylbWntssuMKxAMX2y4QejaWZyxaKV46H4wTU5dzQNw9nggbxZFtJbIL
44togyA9pCIw9Ja7Ji5DESi+JnA/3/ixlv76U1LJuxa8z4E3IJ6e+XHro0JnNpQpiGkisAHzAw9o
7WJHnVRYUHPtrvdQPvFDPUtv0VsgPl5WrHjVDjq3WnAWSrV4xW9C4ZepIpBqJYYUthi8mLru8xfD
cPnuYpZBww2VDlFg9EqXhJz3iFdTdB/sfoM+9keMpZbKGVLCOnlgNn4M+R8J+ETqBLv+J/ECh8Tp
AMEKbAX1CYShENo/I6nimYCN/RB03nTaL0i+Qaz0oOBFD68DG50bTuRIIvam0fEtXgrvVV2QvWlR
TMr7HiVFiC8LR71B4KT21zxzkI0hUnfmwRzeDP0dmb8HxruCeJQsmadzwwk/X/HtR21MB+H7Dega
6fycsW25el1Zk59WWh90mT0UqmowW/5dL8z+GnzjeUVGBb60vpst/81i8Bt19m2rjNLvBgMsPSij
vu8VkRpkthW5qkee+0W/q25C61X+zb95Dyl1bYjUUgDPhUtYds/EOOIMN4dco3SVUtrXFO5jgavh
FjR9sFsDF/31sWVz4WrueDtiNnZankmiKDols6vN3DKPrUoIYzlePgX+uA5DaYJNph+sXgvcbYs4
9BkL29LX4FpFC8r0i58uTg0MS7QMEEbT4EiTT78gF4a94DGQns9uNTO9JI263Bo2BYKkZc5XQ/z3
ULbxN0Mp9/kd/g3qiNN5KeOU9To7PEmtATmh3/huogzNxRBx4/zknUdd+ahU0f0g8n7S2IaEQR0Q
2ZxS6TQ8gABKS2Y2eU9m85PxWp2xdWyO+8HpIack+Q64EHfxy7kaqtggpG2VRUNuhpcW9RwcvKVJ
pqOLdLG5XsW3nglxpPkI9Vc5/CAToz0SVuvwmADIJ4PfeMuC3Wx1pIyFCLpaL+Ks8OZO9EaEsHe6
DsotWCBD9t1OSKlAoGlw/WG59D4gGZokVBfx3cSCDs27iGxsnjCOeALGqk4cvNvJpyw1MrrfXbe4
kwAw1UnsktYS24KOI0vbCZnB3FbyIEqM2H/9/rMGRGe72xElyVnWF7QcBX2Lc66ba/kCjboohQDR
SKvZAlAdejIoOOt3U1lokScWBGUDfRc00lVIJmn2m7C2eusaDjClA+pNYgmDuxFEDnAf/Mnw9MTc
JT9bDgzc4tAPOVe7MteelNyayEmbe97fcc7IEAM4HZe/pEXwkHviCVpeufz4kHRtV9IWRlmN0p6C
rQ5Aek70w9ypFbMsjsz1E+oWrWgUUN1+6NQCZrgkv2sGazKeBve4B3DHo5JmHsFzdwRHhp10yYO3
6HZgDcbm8Y2711SFnKF/5vyMAtK4cAHGyqQhSdMiLorr6UKC2xCsU7G1TqOPU7d7prZcfu2JQhGZ
t2uw8aQiXcVqTGOMQ5VkWSL9q+UfE6r3o9tEkvqedqHaHD1on3U+y2zEOXBWqbDsnmq6FmN0/IMb
Y1xI1NYtmpE19NTGrPZuzoQM3f1EjSWLzf0bVJ5HHYvSDy2q3/ke4mX+/8V/Ef+kdh1JmXbMmnxP
Y3JGTtVRspq6btOo6Pmw1/xe1mEM9+rveHNHnfhuRAY6rMMQgIE6E18aBgz7kzxgan3lbs4Z8Byr
Kf2fAz0eRdmv572DCs17Pc6RdG3HbbVvH1OK0ythhT1jiV73hu1LJO1kqqbFrLE4IAct7K8qZqlo
rV/jyhOB8uuwhmiS8mxQuZDPJaTgCoVHbCyz1X+qnSnszlYHvZmQhb5Bmj8U4RNvUn4ml0NZsYum
WL6SgN7sCzRIT+y9k2HR0FvzbF02Xb+zdhPBreB/BgJLRfvy/btWK6Sl+4W3fO5CHOfo3bNwQ1Ih
gw9F1Qg1th5Cyu7+nLX7GXc4Bim8vZB1rX0qYSxdvL1ITx9egI2Bl0iT/+rXGry2xBteZvXuedeu
ynkr3DDZ+t+ChruR/EWbLG7WAulsxJGEAC8XymDSCAd5huIzwPwSQmP0BJpJyqiNo0CKwzgcXymr
1K0Zukl2Ne+uV0RAlvtv3Ly2lcpgZf49TSemauxixky0wmP0SG2eBdK0nz53sidc/MOvaLYU4lIb
8bD+2ouooxRecMMQrtJVnkL+RKznTkyMGAc5e2EVY790Pvj6OeSH3BXQjOIeArJKJOO9PhJMjAH0
ct/lhp8wudH0D6lPiWXZKbC7zXRbVT1Y9Mrkyn9ojJ2NspCxmmM4hhLQYrrIch2IdQH0lT60jiSU
kB2rfyY0jhzdbif3khaVqPqJYatXQ8dVkRmTj4Rx4adGoQq8lOryJIuJ3K1ldDCOgUKbO6viJdZ6
V55yiZUjPClkyyWP1jEmZ4UdpA+xuWSTEMBdvneMpBctfkjEWNgD0oSy8aTDZP2shRoiAuWlM2/A
f2ORGey2E9yMqmxYIRh5Dd6gVWKzxHIDhY49IA8GOurybekbqxGCk4AHtI4pV7AyMRKpuXaY+GIy
Y/qsw6+8l0/VykROu6xT7DlO6yy3qJ3S7GoUNQr0m9C+jrSbNqhZALOXQ6K5J9Rs8SAGmwZ9QPQc
t96o5XkG9gngT3baZuqnHRU8luR7WVdYGOU979z43JLbbQ8V6cOw+mjxZRscD7Wyrxrm0fzKKwxZ
WrZvdBT9bZul0sto3gzcDUNAluPGKvLHYZDrnIrZw/tdGt4PQSRyoQUTxnmQFVkSZZ9Qgnw2FsZr
Zx92RtJZXIRLGnxufGbyM5AuhMQuhV+Aq7gF4SbclPuNpekF8ox1tVHTy+/VXpu2B7yfdIv0N5K3
8s0Jn1IHVNHzube3G6cVqPnDLooytFidW4Mf1ra14dfnaqSDKbpQv7L+X6A6tMTfdHUAl1FbCJCd
tCSDiCYdOKgVHBdpMvexGBFmEibSauHk0end7PZ2kkuwAlrNsXOGHzaVB64WKOurtew/P0BIn8Bz
Kmp7AUfHrDQvVvfL5Zbu3PbZCBtwPA+bch5bbC324kIGN7Dh0ef9DbnGRG0zWD6H07V7QwFotnll
O4kjvMr1yiQ7gnkcBASEHrM1ZYaAAcrWJ9K9tal8iTerFe33be3w4iTTYwGMM1VdTOw/Y1nxCR7t
5IngTAkatG9Wu9nVZMLJtQFEfPNd+fZPZi10BePKTNIVZ0VQHKl0+9ua8RIKDHsmd0OTUbPpFXdI
BfJjT1P3qdZXcgvsIVdpbwOnRNlKik4ICA2v6/Y7lWbYQAYMdEBmCcUG7SS21czDwvaDeTPEh8el
CL0BpPcOFg7a22kA6loimcXjziJ+uKMhQuMUsMPyNCu5muHVwDyTDYOvgqVhCuNRXtK+XfbLra0Y
DHK5Wtc6hxaHq2C6hYo2TrXnDa6VG4ZsOyXxHS+njW5Gyja7qv2fmWJYeJRv8eOP7pSXSPjaELfY
lSYhdnHGPs7CCayFy2h5xVGmDnVIWwK+E57i8iFekQ2AZeb1ugMRw7CdtzaduoXjua+gIdtB8K0A
VTc2WyPnVjLQD0JY0AgStxqITyHTLRSScS9BPR0jWTLpzXu07hSuQxweSgNg//niJrwPZ4MIsHkg
ixBPpmSWACaATxT2UnGse81+QF04svOcK+wFVvoVq65TBZmhSWYLhqcQ1Xx18h6R/+XaMUh0I23j
ZUxoHb5WOCsAPn9zgw5INAz7UN40ogZYj8dubd8hKrtoOydkyvbzOTR6jbrawhszmjR+3GJJIyMd
wLCyWKYirQhFczRBnGY15fRrUlCTy5DTQ3W4DaWvNkzXT7M/LJ7ov6tpWbQ8jZ/lrY2l5cno3f32
mA2VinLn97HE+MR2Z740aohsZfxtJ2KLhHrlbftX4IWt6YdK7HGngKOF4fiSNHjrjuf7RaTp01de
NXyFN+EYRhx1iDPxuOf1JQrHkYkDQ/D1+L0AdCKuzHb4QAk6FPnQuJZpU/Iz+iAj0OKmKtcZrnsh
rz8wmiij8SuUZ4WG09kKB/8sGaeDDq24IrNP0oU9sW1cA5ap3I5FvbKjvP6KoOFjTWuYC1g7LOtd
B5Ha2fcNE4ZPA/uHKd7j2dWXSEQyk169FwrobckK/1A8npVAiLSBmgr765bVmN2+8XvuPwvowKO9
ooVNVYWauFrlmr9etPSDV7UzW8GpHl1tQAd1iV7M4YtsQH5MxhdLKouKGhsJG6tMphsf8XNiCkyZ
FFJGoANvzeClov0tZo0x3RUj/b+4zadKM3oB7ryOiloxpajfZMlVMT9p0P9ffAObZWzSmWmUOfSV
6SCn4Z3NQFYTueVDbmZBm7Diu02mvbBZrWOAF/6458DMYdk23lz8c/BMQOoO0EG6b0LhscMdgdCK
LOE6QxC6vilHX8Fnfusbt9zO/2MmPCYuDFJ3nackshI/TTSA2hNBEQyA/Q7s+FXDRKolRwSc8/tI
AOAGuPZxMPbUZhSVYN440G2VzRISeI7QzBb8Kjgst4YA7ruel6+BxJStbAOFBwr6IzSaXM75iTMl
PWG7yrTmtzhb5dqIy5cxdriHrOIcuKrAHeL6jT6Ot9jGHA2SDsNOj+TtNR7wZa2v8OjOM5/J2iIO
aH1FxAWDwnDLlwOvELDj7nKmnnlRuVEH2FROi9ysB1Q+GLq+6TBaCwOCu0h54cId83Kih9RcCoLf
z9OKVoWU1fOctlBVQYbzOQU9jyjtXUjr1C9oIfqY3+DJ9F7Jri5pgkQFRoB+s0jONUk7tv8PpB8U
o0tyhJ94THukRW/CSyupCg+3e6k6snxL/RrV4gOyiZkiX3f8bucAPwNdkXFC0VbrjnjtmUCFlP3q
VN/Lawg2rRSRMeA9t+p5mzxFrYtb3f9Qk8Lb+UoPXG9CjaRFJ8YqquaierzdGhTfUG6QayvGxjV3
K03V3OZlWMAnZTvyEeMJViHffuJH5NMpOIXcNqQb5eA/o96bN9rW0rPw4HYhIEw+3jw1tnLjOo78
Bfzz/g10m10Grp8pCf32BKxINgAY+VCslwy1vwQ5Ki3m0hMZUcyiy4Faxxl3GMHANqCfSy1ujzdh
dXdz9VIQFLwgTL/YfFRmvVGL11LSvQskHPuVm0PmS0TKg3p4MpJEi7EOHctC2heMnT5M2s8CJUla
g0cYr7Xi5w1HzPf3Yf9DKKLiZzn4VvZG77ZbqysydRVcTqfdX3kpwniYnznmWmDLT3c/6c13ehw/
R2trkJjNUxIcmUoKFFH2UIocyeiXfOmh+AnUiedAmfpXgW4NCxXZ5Ezky04pFmAjmJjLm7mdMFJM
+SSnf4ES/eThdwq9To9D/n7jQExdhAEPQgCZatgj1yuaSOA7K0g6sRVhGEuJOrpIDIyYHpMSgEtX
vqsCOZQ3Gyb+Zl7LYIya/lDmn51WS4HgCkzfCUkJFO3xPQidnXHWKvQcKWWLGLaZ/arbneUxZiRK
EHnNMqSMZYsgkoeqZXwC7js93nz+We1hNJIOntDf7Ba7NCGkZpZjb1X82b8bQFIlUz2FteMKSxcZ
0GZguzfN00kTinYTKB8NNmYlK4AS0xRmoSECVmtWIVBJeHgicvhH1l61z9/jgu6KYHeFSdCNyg/D
Pm8hdVTYIjzPgQWdzjRDbLMGqH7t/lu+XOcHqW3xnNjETAPWmRFNuOJ46B3wvk4apCMafRBAHy/3
hhqyOUVV71Y/LYN4gtJeIrjMcWyndtwtSG1YmCB8vGeprRDCbarLdl6XI3MwDnZQHhVf0A+627k4
TxixME4/P9ICH6vLKFxcESo5/XSUFcGnWCa6qsBTiR5TXjFnRbXfwhFH3CYgGukZ3wdRtHDI3NIv
oqz2iXmfjB9ZFMLyfHEkV3STcU6Ww7LKjj7CE4DSUsVk3Mr/c9eXFd5+dKnlo+d80nRkEY7b5bhN
ppa5D4EssgcJjU4Ldkq2mv8Z6YEltmEjQlp4AtiVD6jslBpysl6Cz9gWsve9DaQUduPAs7vSfJ9Y
SssCuQQ1RsySCPj4yUW5g1frQtwRgch9GFeqr9qZftxVuPP5Mfo2ND7JUo9vWnsSzC55BCV1p32C
AXTHnpcdtEfb/lon2lvT8TlOwMdlssbRrpY88Wcy84MS+cmyzopyurHRTe2u1N85ySeUw9T1YZc1
mEGBLwVLNhLoIW2Gsm6Nxr+QofIGsOZuHpMD/W7GThU5OmdRF9VMhg912MVxxFJX3Wh3D5K7+GnF
WK8qSxk46ot3ds4uLHBkVxUaJUyPHseLl3s9q5VLXvm5T1SkMViX7C4N22zL+oY2udQGJrZ2mDF1
osycfbTfBxIXOXduzKREILIOdYNWpq9EPxEtcw0fvF1AOQgHaGbqltEO6CB1yRb6qQBaqhtgFB9v
bGbjB6fTn0vVSHeXqKJJKXcevDp4pRw1zoT6LxeTdYWIq2pRWi9gK3Da+Tqt4oo5Y/srjRbDcvGA
R6ne+YSTsRYotB28beBEg8I3SI7lFu5HWxfeqTpoAYWvXrGg4UqsN12qe1XI/dU+Qs75sRbKIPOv
a7ZbT1fU9qdAMUj41VI1DoVys2Zh4EJIYZ6Nd30YMj76NleRq+G1/nl7xQSVqAPOrv62ZGxFDYkw
tRLTqnpd0sMzyxxOej6MQeIt4qMbYVdBTCBGbmsxgI3PVTs1HQK9jbb2nagf53cDjWeMQ3RHxRaR
tzYrX5ceEiEQjNsiW6GGNnesu8t0XfHNAxDfayVnFkN9jTnWPpVYOe4yT7gZRlCMTdnoX92gXyjG
ON/N6Bg8sTrFNKkalYttYfHVbjI5WChEb5yp3u67/Q94s4/cdb26BR97AeCef7lFyY/pD2opqyVe
xpCB9Ofl3YHyyllrWd7blDA1hT5O5BDfEZlm1Ln2zbfsMASMreJ2A+z64eeWt7WqP2qxqMmtSSTo
LvoOpKQFePUns1vmw4EsKbpg4r7Va+LCdCywk+QGTyu9RDkmaKVNDA+Fsf2ukgLI7WNG64TYCp7+
KBCI4pgTN3970DyhE668ESqBN1eJ/ymQYsaQ/pdVkUE1Wx/Gl6/agBHiDtc2E7UfMGqaOXrv14xh
DH15Djh6HJTpBeAkI4O8e+LJpN+ScRdTojOPBSJRQWV9K4dm3HnOBYrCnAPesWoS5gUMPWw92Nrv
mhCN4Wf0Fx+05++2fJAgTAOjLKyHhjOLC8FBo3AUv+K1uyIgGk0gIzeKE+Rc1HQDqlL0/jABkEJM
K0abimnD5NyiZeDHjoghJLh29Xwpndp5bIipnB9F6L08oFOsVDdDWt60O8R97nGDWhCuZmjInSBy
m5LOEU34Ja98jiCHm19NPt5iOpjzmY9QcvaBTbzhATaksXloIAE3ea/W9SZRzOkUbRgz1/EyRuL1
OryUPBOqbNqCG68sR9fxaEAbG1soVX9O9Ka9mHiEni8iG1cYRiU5wvSSkvO02/P2khyrDPSn9v4O
B2Vxvhc2Hu3OeT8b1WEz67V0TPWpKjxzpxYdww47DKzqBfe5DtMb4sqPFwQcg4BDfG7kB7Vp/uMc
vdOAaBIZMYibx7Yj6K9N2GhuuAiJQIzbVyvCenUU562ssjHTzszDhv+BQ4E/mKb6irJzFq8wsUiL
ZCEOvxRhzISDMQ3ku8hXSsF3AKlnKFZ4kyHbyTvMvNBKxs76uIZqm9PBVqZBB9qs1N998Fwaitmv
tmJFb9y+tc1sefncW+PWcUKTW9TCQF5PX5eCW37BsTGaMhwbUaNZtB18pbH2eLeJIOfgBfnwdDxS
EWp30DqgCkwiwcdHSOmnZSxyBRv0xPY8BlZI+j4nrPij4Hw2ZGxPsr/BEXAlsCX/QWryESIBPQjx
WDVSFd2yDbfj4h/RWO3FdFcUQP5OpjjKxer+wwP69nGOEt9KKr68ZNE1EKjYn0G2YmYROl/bcvb9
Kfdsx9aJlOYxutifua6E2Z4U1DKb4ELgvYinnz+19h57D/ctFqcuYfAWAe8/qyOArrrLi/Srl6rx
4f0PzXFj9ASgjLtq60t1eH80OeoVnjE7XcmtjJU0aUO7wx4kD1bFGPqkhCKMFLNjQJW2+uVUkYjv
3Sil8jIT1bo3Np1wQkex4N7Td4llZdIVQjRIXqqd+JHeUEe9+pkhvNLfz+bw1f8MKlOcb3XzUrv0
7JhpYx93zcG3CNEnNAXI5SRqQLOureSoKL1l2JjwQjftgfNUhvyOOnsoQXy35AXTcwDEGmSAIMry
ajAldI7uDtkcFNsRpdBUM6CzCRyKM4mv3lXhAtRVIsj78U5DQJRdtPRoL1jPK35dannTXQh54nXC
wxuqD8Gt+Bw9yWK8dP9Q2LOm7WQHjBC3ZFzff3XyBcPV6VwJQVxPJDMQF8VrAU2dMvPZY+Vi+I55
pn41wADpJoGLQVtoOh9VtbNVSmJLKe65yFKTFnZzoMy2LnanAIZoLOpjryj/TyL7Go1o4JRBpe/K
FEp47dqQ8Slqr7Nzo6fSEcfO+VEY2IjSJcXUSlqhJpGdWfMIP0rb8oA806CZ/bpzfYcOKU5q5s0S
ULfHKHyX3IVl7x44ETZ4FAOaykm2zJVmGX0tMC7RBA8T/lJ8ox8RBI1582S6paSirS2qnPrj2uOy
zt/VitbKKh/9jLGYzCjCE/8gExaGNB3u9Cg1UuO25h4H990gB37JWeJlDQV/CB8XDuuKW/rF1IMC
08QUBmDIqGFUmajFGJUarY67hN7rjp1LZMvgV+xi9wL/iZ+CIjb4W3lqDIbIll+urX8+RjW26rHI
o2hkU4Lhz1JUj7N04NaZ56rMBTtwTl7zB8+Iiyzojh1cDL3FBe/UwqBJMpbzyl7oBk5V2SPZasPC
lSOyS3nPf16vcRmtmZQa6QQQjF87ibemySEMQv/yJts0CFJrJWmpohNTWwvBwP0pSi3Pg/ifgUkz
oSwR1VbPGysc6G2jojfSKb2ryIJNmss/2O+F7lA+tZJlxHar8OxOYq3UXQKE4yi7xfo6LSCEJsQv
al3+5diWL3B55KhBoBbTkCAIewpWQ9XdBb5mlj0rUrk/xv6AQC2fmGuv0cyIbrroSez6NYmCoRM1
2DsrB1tDmbnj319skMX7b1gOtSggxzFCLFgjddmc//glcMbEgEX6coW3v5VLgzoPMQ2DddxqFf38
xIbdpxMVU2jYPjNN05ZhDBaq41OBfEDBungkDZJDKa+pSyKKSbmImUXn/doROrQBmRlGZ/wm3Y1Y
2bcp6gdBhTRCqvZGxWyUuvurL6X/n4wnopboCUizy8XJW7qUt/tksMI6M+CAtnzH4yRXux/ARIAf
azCmbskRDKt6mtvx6SZMNxbe3YnCQHd+MdMUhPqyfZHcYijnQAuamhrg5OdvysrWEQfeUK/PyIgJ
VHppuQNjZYA0OEAPi/MdtcSSmM8jfCAL7KWbPT4OIc5QtHmhyvs+/0hakwL5SYMTKy7QCuCo6C9i
YvOVcO3V0jELUi+ybfjwsmoa/USShQVCEnAI0wjngwXl2Kkre0/6uASTA/wr2Vcvy9R/HPEXicU4
cdNKRzMxxoPslUS4ahkfFtxi8TUm6L9jlFCs6JBzDHuN/qthipM9uOKnOn3PkJqle3oa3qhl2P7h
75K335SfBMDdoq8U0v4liw7LQKp6AS4CqIqzzfLVG0EIbg9Gcx60TLTkAARxdI0Wx3KHM5by4Eli
1tVXk0oR8PSrdH8bfOXZkFLlBe3z9dbFBdN6I0NwVSra9iv3ouxR4J8PEj3nq1YQN7p0+L2lxNyE
/fMiyS1kQifXQKVxdF51CpU8RYWdVl1te69YCahwUZcjWAS0nebi/zcIqCAVIN/x1gK1SPn8YYDW
UkSpuARUDXaXyyGLNMYCCd4zBgpDpjDwF6NBCktzUPbTRnE20MC+JA65lfpTEU2NlScND2DP3zs6
ltbbVcnPmAk4wTmczNGEy2ksQbKEpFAQtq9DFqOeu468EeAM2mb887e4+T8XNstm9m4zcg3h6mDE
GbB/X1iSQW69ZXV1jem08zCYigGqxKxGF1qyknS0gCYzW6Kc4VaHLuGAIpPDkdz3LV4GLB+doeHo
7z2yXdzL/jJthgCZAlXVs8t9SDBxgkm5KDTHTW9Be13tkGdzLgeJVg1dUoX5Eb+7HkgLyfWLP95T
OokH+zRvfzTO3Xg3RfvJlzm29l1PYH9Belv6lVGartIG/qoqXu8CRmAOj+4ioF2QwU6moHuj2/wC
67NL/cDt8OKVJ1k6ScqDaqysK75q9hJ865d7ZDxk19zb/zxK0bjPh9h6kSpQQcLhHsdU7wsdGiRI
lxkX35Locs6aFoDQjOAdmEuNCQHnuOrX7fHhIdrElnyK22PQDtYRyMpNaKs6NKNnR6YliL0ouAC7
TO6cMveTI7pPZsyH7c+TRGMo8YceJfisOAG2T5gf4iZkJU2pHNGWGlkbsc+G9sWVU/EZI2UBd+hJ
k+OvHs/KiFTmv7Iw0xLVHt4IM7Zs7pqvjO+DM/HJAvAjKSeSPl3faTiY5QvwtgjjMtCOQb/Mie/l
k5NNTMIlfBUkn5WaBynhWSHpGFse662c/yLtn87kCESKaJLqAmKeqHaRx4FaSkSOCB0xi7+K0/4t
wybM6ZSXvwy4N72bJ5VrQmMppK7n7/7j1BtfLaDZlzrFZFy3/Wdht8pw75mlTke6nOeVcuf9Tlkw
hL08yUp3fJARgsxFKIAdkB/5mFcqe5wupohOSt8O+SdhmYDNzVKAuakKmKRQrNCtCMfK4ougn+Ea
7e3KN0gXfKowmBtWYH5FNePca4p2APiyrq2ryzpKGPK6Rh3q1Km/b4TXM/gKkble9Y5qChKl6YbO
kdaoSINXvbmUXj6wVi6b/Wp1215fhJBd7GtM9/4uYWTbWlnmOkOSbRHpmHwBcTJpCsu2IwTuNSYm
JQkoI60KIsHWksGIE68IpiwO1rcEkyJPCH5NnRSD+78LSXwcZTtbWtXBMgWSwXMnDz7jXvFB1jlO
UtiC/5SuSqzrAHDH9Nzwvyh7xROh1rm+y5A50o+9D7Wnuvz0t8Rgr6kdQ8ks1DlbpkKtWVyOISqW
U1wnRGH9N4kXO8M6Uxg7dkHsn73rXMv1mNIfJfnZtI4UYaeSH7L+F4+Lq4mv451ofLbmeAyTbD2M
WLFuv/fCA0yQ93zakW5uiju7Dx+6VyXmtTy+lEhvyWaP1VpjG8qe7ke1xeZVITDpvgrMDtvEvBLW
WW7k2EwRaXLUU0QAymeeDEGtc5qlU7gGQPm1K7QeoFDo5agG10quU42fkgTwOuK8CZQHYf6+oNAB
9pzVz0j0ez1hWsIfmSoO5oq+pdRVTqNlRTaDBfKqYBj3Z7aAeoVXLnnB6CxPBTjXzGsq501Flhby
sUSE45uDUCW1SoO9uqSgappHq7MWyjRfMUOGKAONSUBsfI9e99Gy2mXxJaxrEFHA+cvp6NsO3nXQ
5jsMBywi7GEi8cwHum0ip+bhSMFZ77G+J7qlKDCETo7JM9EueKucB1pIuyOEcKPxwpZY1jHNVBnz
t9HgwgovBP+VS6JLOpXsRBjNJnGcu9Pz0AncgNB4tuSiBjUiSwvkTExsNghj4wkH9uLG7EawiLHe
lEnAMZhjbTlMdnTfys5ElDty+SqSB+MR5ucn1v8uFIF8Hf9ExZCDsNTJ59xFSI+5n5CHeKazzZRp
+pudHGa54UNjsKV0vXNHFGfuORLNi2GXy0vQadZQu3NKcO1NpdZnnpJtM4gbjj6su9uguUtRVkoE
+YgGRW7iMBmEwI2la1btk81ySMCDYJMfoz9WuqX6yj1y8OEYEoL9T0043tVnLG8WsLbaWvLqa6bw
Q6LSNGuVM1y7UZ6Ur8NYdURZ7AveJAUd+KxMdl5oV7QG3B0eNCzLm+nFFPzNPhq5e2WEeVX8rHOG
jUZvW9XtDkHgbBiT1s8E4mxzikR/gBXbm+qFh1uIVXbGe6G9RcfGy/pMQqmv9XkXpI4pNml+T9o+
o4CLAkCJSjo+XYdeRLtIaYXCO68oL2W9BVFrFoZV0ECJkQ/IFBoHX83FhkQY9eP8hiy6UrsBl2jT
ve/U89OlkWZEQYMqb9Y0f22RT31ULOIqLL8Jf/e80qtTz4uTudCJJR0paJBKyPxmy6V8aWY6Aqsz
6PYsegKS4K+XcyvTiTh9qt4uXWJ80T3eBe4E+O3x1anm7wd06Gk8+QTR1s67uprSqiqXDe81eSIW
872xSq3giRGYGTEQ8/ZmRREhUhF9kENu94Q9AqJ/n+9QrtPWzMbHvPX6FC4AOb0yPL6KEUvpm3YX
FoDKGWUBOgjs2JILy5EVQzrJY0KBuH8AJ7Vj+ZkKjTkFOUCyVZkmkxBvZ2noei7Tbh2g7DAVkf2b
5JTvaHWzROf7zOWruJ7rQVAQi9Rzl95nQj734V0TBXV2eeAPbOwNI/S6ZrDe6d1KAbEHctlQBiEp
PVUPJK21pJ575KcKSj9QWBy7q8I0KrY+nWO5lhtT8VrXWN1lAaoVS/uEBEz5e7a30VpCGITyGo9s
qAy3WjjMiZhR0YmoBFOg4PkO8WUQtrInNcjFKrMSUl5rTpGHR8eWm8bSQ4+jzowJyx/9IV6Qro2u
s1UVONshVhBGlLiGdFfw4un4g+CFC9WAhV2f+aYdmm1KJL8VvJaPtLeYs6kILNxXgQNeZpT+JBd/
s+MtfNvdh1Pp86rNTfXBW/dF3KQGHtk+ZPAxCjPpKWcbVnW11ZyRU/YdWvIlUiLjmLs+CC46a/Or
/ujM41l7pdo3aZxRynLqPhoFk/hm1XO+zsmM1EdI72MGjM07cyK50xNWznNvGqLrwBVn5xsA0Tuq
vwxOblnEvqAP2Qv/oVtCAcRHyXgxKtU1e0zZTJTfLewXLAsZntt6K3oIbLKtfO2VUYUgO+s+SLl+
45xtoYBKqgvX8GxuIFwb6vkPG1vSRSJAcfTmqthwh/x2005j4/VLcmdgx+eFPlM3+4/+i4WYzd4R
ggtJhy8ZNxZNXIPv/i0kGlv6vIzWK9S83w5Umf9UUNoYRFsixhBuGVJlg8wii4GINZXxLfejw1Hn
7vg6g1I5uIT8X9paoB7GFcltQgSH+5B5DQ9Kfi9DiBBqhBN6Ysx9PktQvhe3TFqtK1cVaFs5mPLv
UwBzstA4Yn43IJZjmGy+FwM8iRmOwOD+sX0jMnAqvy+RyJyp7g+aUQNPJv2N1MQG6NHDzym8mVvG
OC8WSGPmInEEaAdpAWmYu8nuipkVeUPg8AkLdhFrAZjfBbG/YaYZsYthTtXAxzMVc4fvCON3OWUO
89X26CqPvf4mG2KyvuYUgyYGr9Ainyxi2vOuMSu5DU6bN3iCOxvCWS52L8UxOdI0w7vsU2IxKQkk
7zg4GOpAt4qUsFI540Qq3GjfjLI0tZN9iNmLzlg1GA2Oa8hnUEwg/RHPSBglq7Xb0TGCikzoOA4/
99sHBsxsRIn0J7aYwREF4LHWtmzkL18yyq57rKxgx+Pd6G6v8pLG9WpIVTtm6b0oLmTRs7aPI+nV
F3rt/iptrNrNYT/FW85olVZFjbTOAC9AJhslscZ35/Umg04Pl9bdlVbN3ma2mLY1BLrXLUjcKfF2
8ZGks1RNGPmaAG23NfmRGIImPffzFRNtoJvSyDqtFyIX7NI6xqRU4UDdeFssYFrTxVEHq4N6BDtv
8qKZAKMYaVwxDskhtWace737u+/25NEwa+etn7liTSqeKFdXnnTgJgj9DcsSQj1Ws3weQbsZEoZj
FFW6+wdUEp6Nz3rkjAys/Jx7hDVHGHPmDJVlpoCvTHKzVLZ+yKpHDSz1gV2cMlyGtDlF/XNpZ6Xt
36Usn12w560zFDvCtm4/8qKRPoYCmv/bCk/8iXX+QsuTPfb4hPNWf//N5bolNOdiX168uKKS6aZi
vEVzL5U5ewAvYXGnH0iDcTKvq9mCLKIs+rXXGboaRsCVFF+jP91ezjL20avmKyw/jMxztWkogXAM
wyCZyiJYb2uFFl2r1xjQliA/yn7iMIVKSPWLWipwZBk5cYoioZOEelOg7uPMx+M95ouYRFO46x9V
swXFVSCVF3qjRBmyulSXt7cB8zr4JF7LgNoo/J4PFsL6qn7dqyTQJkuV+DNFCtnJaf8R/g/Hr/RM
SBKzIeqmzEI0R8LFQnYS8L1XJtHqVAZiUeemll82TwsHRRXa/VpDiylBQvud2WL+ngDG5PaoyJQ5
as/HFU2uzJes8I1nX+S3RDQUNY01Rpt09aN0yrvuD0ztR92WrkUMl94zuf9QVEeTK3pSIZdDhrnN
orB57GWebgrnOOEqOyDiz0iV0HdlDqVIxsP1iHCwoJoFNt5dXwMr+xsPgzZgm41WQ9UcSjaG9ezQ
GKM5ssmdRVFOLMwZL1PaBia8FVK7cac7lP7+rsQU0/1xL8u3B7SvVusEeKkVtjjyfbmFXtzMDrRL
UhSuoKf97GB0zbYtvZddKN2lpsca2DGMWi5inJqPu+OZTkCompYMOzi4YSI9SO0WyOIKf1oFDqHy
naRD88I2BtVGhHaumJyI8o/Mwejppc4VuzpyLde9JjF0fjWVCNCArr0SyPqNaum78WZvi0e6wmn8
n3O1dKpb5RSWIQq1FbTqlRq61clY0iJOAr1Y/1zq5g0YAxUL3lkgO5tmZsfnJl4LOnvBZfhTQRU6
KQBfSYX69C7hsCT6DGnhCCrDrI9G4ngzBKVg1ipL9ivQ4XHDSVoFaiZHQ4wsNOuJXYKQzcCFxtAW
viZaerVuYsUNi7RJsAblIQW55vIae73C+B+CB4LDRdyorC4rrJ6UcqS6J1RWlqNCJnrsHRkcJfar
h3FfDdmeVEp2IldkROAvp0G2xSlThYDHBuZP6PlXTWqd8rt5c8Xw4sIz0cxzchkDSM8o3nQFcyzS
uH+3OfY7ILbIeaa5b3U96TSjX7tISSImC0duFCaDfLCZ8qcxmdgFABccTcjtpU5zpT7WTOmG3wfe
t1MnhMQY5bljDU2X3aLnTS5XXqi9G/VMFtCS901fTl0IlUrsDYV2ERKNkApy2ntsbyeGfPgfKzlD
GN+oeY7lf/+SBhSrHR+3POANrnpxY5zvagc2HGgovkYdh8/wqJDelwRt14hLDJQTYk72isTiVWcr
VQwK62AlHtWR5CH3NAMT2Nu3PPXAQf1Y30GBgRJ5oKRAN5fMTXjOIWZLaDCpFzmPla0UAwI43C+M
M89iutvea0ySQq777r7TJXC99+Sbl/JS4Z6Umwvmk90fTpwjHUIooTdAmuJ4INJJQAVlsvP5vSYf
s32Ojxr9gH0fUqGp1OD+YjqmKJkuZLjAejkY6mnCsfdO1dt9ImeTrFVMy2J046Nq1eCC/jfTNG9F
aCqL2dOzO0vHbdoeEuK8Sd185aBJfi4OW+fQ4cm/4bBOLXU27pXvrGYXKbnQujcnn8FOstuIKJS/
TeOTZfSkxul1i/975xe7Q620RhHz6kccZYxT5fKP5hufYUoR7qPMnjQDIOd6G5Z9QNdvAG0GT1J6
wThIspltyFMJnvsnJJd6zocs7uwRjMPf466sT4Re+163DdnxpcxdykQGZFsNfLPRTIhkrPEDmxur
qjmv5mVlwuMQi0V2NjjM+ZpleJHwzZF0OyOiuh0wLdzd57la8eNGIfkRIxrSv2iHWW5BN0H4iGcX
9f8KL1I7Im4djZG1wo/Nuv0LJowvUOGk3cuFIhr2eFTf8nQgeaCUS0k7UVfnx5bspRRWnFtIKQlL
8zt6aX1VgZX3LHa3KsAvYx4fvid/t0Z0nm4+pdSnxVnPA2MhHpX25VppbtnPmRQDQWcwfV3LtZga
C4aK2w8/oJC89uMqcevtg3ImsO4DbLJS8JzmrVhJLwZaZIwG1q2F/OaddA2+M+mcfEi6B8fu/S13
u+LeEX5KLLyEMgIu1rVm3qk2SqehmBZ8UdmFAA3TdWboD71Cne5E+LlbG1gAFen0eWUoIPjFPiV/
BkLAgzI8VsWpmSb0iKrMqVFUyhutAJh260NkNER2+6DBvh0VyWXu1o6kLo0Uuydf/cfRF+j7F/Op
W/BomLVJ/De0sOujyn3oCbwvae8wTdSXuviizCT7J8PTm2eqAXrx7n6VQ3AIcuNyFCulMUa981JA
wxpNOd8iuIB94Lp9U8oU4lNoGsCoPYVh+Mr4/ThYIqSUiRInoEg80Ah2cg+PXAffqlQflITxGXHc
oWEhf4i68KBZVuDdGtq30LVV9YRn77SqkoKYN6LYRsxtBZG7ilXwHxx3XmP2BDA09op17iAR72Gz
9rkhxQKl7YUY4k598KIn05gLhxqkKxiTkQUpnYjQOB3E99C88+CGezVTURkev7WJ9eJEsNB2mr+z
Gx27glu/Z42ueZ1Foo1TftS540S9+4Ds3rqOWahO2rFiA83YzzISEkPYZX4JIYc1QTYeXDypN4NC
azViMm7V9+sZVJDkak1w6AtnqdxtEdLxK4tbwh+Nd0RBH1eaTA24DNtORkWh276TiONik/EoiNV9
rCjR7ZobcaUfBiXLYZHzoMR2HEa/14fRJo+MQftF4afjkhQYOVPZ+ofglVlTb16rWTyK+ns/y+pO
ifo6r6JcfLrEqVimgPxjnydikI1HqQ2ct9BuP8VLjHu7FYxo3PfI9Tr7ISaSTIydFPUJAKYne1/m
4dAIkjubqzg6nUcYYO5FghcsyaMNW+EA5KOJhJ02q0Q7xCUc4QGGh1RPLhB+V/FrwF8hk3TBfHG4
gKD/CrZ/5bDGbca0HZ5KN22yWg1tORdpjh8z0fLkKxeuCjLshTMX77k6zXl2ApfBGT0AotdrPJaS
PTN9IDcBfbodwePneQcxE7AtkjjDng1d3m7cuspfwoDuOtws1KhosrtztYbsAXGg94mgm28OwO+Z
VLBrVhBaW7XhZxIOGsmDICNToY6xggrBayTi76LvcGzqz1EMe3RWCgcl4WbY62EyrITwI3kE7vag
+W+0tvHDlV+2qdXiunELFuWXFBhCxVepADr2zNfxUzJvlAv2kncbttcM4tnCN2/0Xq+YjzGdLraA
wccBQ9PJIn1M0aBc0taLB7Nj+FDuIKrjc+MHxbrDb0Ko9b/SevkAq7frcNuqxD1nVS+2jjecjC+r
0iSF5oVaHPJ7LZdL444pgSg4uCnazdp8HKD75iCsNQyi5XPfjIqB/+02Deh9bIk+pWYv3n7IORAA
+1PRnibu5RXj/ra8wTFvIAbf+dFa+JydwZcXiUfcevcn3V3SW2VNGQkXtXjB3bRGTFlLG02pTwWY
I1pSH9/z5tR5Fj2c0OpM8YMydnvo4fLYc1cd9FTS4Zu6JdbkXTQdl1AdMB1nSriVfPWRZPG71DL3
J1ndXfDGXT9qTKdRgiJO3eanaF9xOKF5EmyCKMnkrEY0b2g8F6+uJy7hf5UL4wHKmTVF3RUWq7Zk
k0AAokpS6Uy3QpwxkfWfFzNkkLQcmTctJlTRv42C0yK/V2W8mqT7LepOpHX23Nj4YOgvzF/rZawP
n/Oy4AvYENB70tZNPCVA+OzHCrgkOBGzXG/o5RqmVuuAGO/l+1eCYU8oagZjBfHQoLeYAa1bRRrp
8IXM1aGsBa9NsaMhIKkM88lGrQ7HsU2oQvNoNqNpu8NwLQc+a1Eez50bqMnpkTZcykjYRecLWh64
4Zo60IHiHnVFwPHKe8Mqchs88T8ZOdn7KdnRi0s6J33NV7moiJEasS7kiTybUL5xpqTGFt2lwEXm
KybJThAyzXQpxjY3auC+cK673k7r7jQlWCWuzWmozmje8vynLeBWckWcqe/IA/eb1l0iUKT9OxJj
bLdRk9AauRd2PFNfxrLmSn4LTTzg49fkBYcnmzHCtJdcdH1UzvJssYBbOPxtJg+8ThdgZ/FfPvrR
X9t4KOnaEsM6d7M33widvNcQojfzQYESSf783W0+GiNdjoK/2zaq13VZmTgpdYao80pTIbk/jlDT
Sg9Tizprc84yUFwfkztuAqoqCfn+g2F9jUSg0NiKQVbi8HS5QszAGyEpd420Z7QnOtDHL8+BBmVf
2tTbsXVRk1ttxiD8S0QfQNRcJO3tKpW9cvGY0L/0pa5uPP83rJi5UWoKI+ZZkkW/tDELdYhxmXn2
GD/BaITzfpSmycYW7bEnkDtL332hE3np46SZssCeGng8gOtlmHdqNyqBvfEzqsLPpEqMtAjjKCAW
yff3fypJlQuY1kachkGO9LVpU0BmigHjrx5iw+u411L9RH1q8XQ3XtAXNOMr7LHtG8l6hQYuzvFh
r0P8GmiWCj6Ya9s0TykNyiXClFbgbUeX2lOuZ1Ej2he2G5oSBicRYsvC/smunxfgjobleim50gBr
IS5RF/x2aU6j6vLId/o6wy/bAcOb6Yd4DxVSzehTRokl2BAYlot8/aW+LfuwymK2MpW0kiXcDmKi
q52Iw+AVR7J+aADoXcsWCQ5gnSOem5WLl3oKDt2tHVjtTG5xsJ88Pn6jgtldGYL2vCZrDekOiU6X
j+u4ZJnSpIesqVK3eCmzg+jl8ljGgT2ZMWcIgTeTWA0W7RJnkW3tUZvDjvEOLtYVwAXMyAi5w6Uy
Q3VeqDm28FfsvDBAedUIomtAkkTQnoW5DzssBJZNUNXob7SMw35XgWfWxZrQuB73kolemUSRnim0
xGHLz6PQHMuKyw1vZ4Gk+b+G5vUfQgogYcTGwaw/CXSeqKXC6sC0rI1Gkg7Sayrj8nNVjq3tlFU5
GnmYCAxsnN4HUPvBsLWCYNMclcW953SFyCDEadIaTC2dbd9g74MdJEBODQu3Qnwsl+NhQKijhoSD
CJPbLGaY7rqu2aQ09JSi5+cPkmAvYD/JjlQMEsEdaoRtNlZIs9KQJGHP0HvBY0P7jt0SznkBWkrQ
ogDahF3ScxNI8KLHns/vkbzQro09Q6YC8dXdyJ187e9ZnVqOyWJbr38TJq5vAVTk9AeDVY+q5mWx
UgfuAdV705Wi3jV5FcG0hVzUt4y6z5fgesi4MRw+K54wBVKITFvdu2PAyxAno7Jett18o/gZGmlH
aTXuLMYeuUaEmD9tLZ8Z3edX6dkXVXwQigvPdEeyrL/hfchn+178Qes4BgbKCtGhRyv2yxYuvrZZ
0G30CLBnJDCWJ3/m+DdxTD2ZF2wRxKJrCWnjglrsmFVxt235ubaOQxXRujWDwEOntEpGyBTwYeH9
bpm1PR3MrhWrcWtoQIS73cQLkl8npiLDLFqmXUZ2jxuPIRGZl/tB5ADZbUWVfRNAq8Evu1IwdFEA
ghmXhpre12bGT4mWmExQnDtpfsQLsuJ0ZCK2TIiJrTlci7zoSYwjpenx4rwwoOUr8/8EMNieWMGm
1Fl+fwAzpbmZaVsaOd4dGRLAqusQSVThNbns6S6qtiIdIMfBcgetvmktqQWODgBvvie7DJIhg7Xf
SWBxQXiwYFzoddma1yp22RmS3S2n/je8+A+uYcoOiwaYcCme0Z+Ut5LWFVZeiyxM7Y3pTlVUbbnW
pbegDfMGXnQcP57C/89xlDmQ5JfHc08muSFGJ6mwi0n8yYytTHWW7uZQpbOvn0BqlhvXBGKuuqpp
4BNUcbIvfeQriZqVuXNQXTnTaDFs1mPHIO1dp7WI56DCyZszPmDxnVpRmdjR0Q2wEgkJ878Oc5lQ
ifZe4AvLz/aGzhe8drD+vbFkYqt21fxDh+ThMkG+rcdJK/K4woYOm2cEm4CqIT76nZ3tJOyrCyZL
tWwTRddXYTBUj6LTWKgZTgYPymgyvbIRErxxvJxLlqnWkSRAGFV/Z9FLW9ZfCiQVCeU3nyzmI4Ly
tVGr7FlwIsn4gGhO3wpCShdSzojbg8yQp9dRIxT75ACjJ94oRVFFpelNpBrO7VIz6btse0DOyxii
GqknssyNIPyFdIHGXRci6nkks/XDPQYGUyc3EIy7P5Gwp8i51ZtI0ljEcvM9mospOJRRf6+qTCIr
+yhnlzaKJ8nThUjKH+G5H+u/3+3c0U7ljBCE3yP6pgKaEEMTFAMw0bClPq2SIv4oopwyxSfFVocP
Wpri8HhPvHXDOirOsUq8oeEFfDS5WFNcexzTJ8eAz53HjaqSivbxdSEK/ASL+qM9SGKAO76c9UZU
ypKojw/ob4S5unRTSFby7/WO26C5D7ZVZWAKZVdWZPCNFXgNCOuc6I1RYVXZ4Fi4/eCbtso6m9e+
7qxJgzsZlu+EJTB/ThXOncasA79UC1gIDVZ1dUJJOLCH6iSyp05vY61rPx1h+UvCZVfcuioVVDiQ
/A3pfVTxJ9j498RarcBodZLZ7G/8bTRssdZ40fEreaXXP86SZ1/oZr4XCbwWjwmfjgIYDpM1S7Vt
wqcqHqMDyp6vhHOcK4811019/zX9R99Ds5GmJTbNfSlhQ3jsAVgU/PfD7WUyk0ZCrMbywUtzWkFX
i4WdvcVDXdwyb5nGLgZ3MghIjWKzxpTXLLCWVi2+fdLGXD20b7dPoD/igIbzb3rTVa3+fsalY+dS
zl0vWS7qCAbe9h49jsxGBNWObTC6qTiliKiFOb3J0PyKGD8i0jSAqQOWnDLffPZ0oNBbBZuig+to
LEPiVcNPm4eXjSpB4aml7PhVKb2PEZSDP6cwrmasnr2P0cQQKeY/k0Sd05ADeBy1p2fJhtW2MGUu
0JrnhZsvKsxD6FxX1MlcOnmWYie7AFxATqbWfpcx7PDZf+GpoKghOQo3aL8i0CSL5A2mpg7WTgfM
qx9RAzOD2gF+7mHtgf05k+35QYm7ns5xs+DjmJ9wkP0NSlrXMadbpfFYtdFLnJncOHLFMcnGLOWf
SO4AogGfUpgbEKa5ub7W2KygM483XVM7WwDg2vd8ihM72fyBECAqY03y30wNYPf1nYEu8ukbdAE5
shWoHgvu8FP0P7boucqW4kjbOkuZ4X2bBZPkFndQlUNCjyZuBo/+40AZXJ3Xb6C6NPLwMmo4BEVA
iXrCKYuRnGYd1lCAQiTIcguDeihgySo1Qw0bbwxh8+9jdk5GWdxnMDuk1mw0S/J31rCAOw3leswX
fNjCEcgroVxLKbHT40VUXoHhNIED4+Yaro+dPZ+DoawE9t+Iv5CvQCrVFn11IGjGpHYw/ITcfsHf
OPaBIurXzdAJToyGd4tUKTCdU8MpHYJuJvXdOErYnKkI4LEf8O+cjc2Rhn52NI6Exb3xPpV1qBHa
6qkCFxkJQ64zVfV7CoUi432Q2gaQYxpsF9yyFIwb0v5uDZUA4cRHdoN2RwnbxrY/UiJnLguzuYu1
7vBKeea+tFcUD7tjAQEd0TSwcI3LIqKaW5KBQ/j8pf+1FZR5Ishfx48OhvxpTu0v7EcR93ssVG7d
kcRGDZkh3AQMGm58eu5lLuqg5tw4+13oi+uqER4DiPRpcHZ4Cn44LQb0pKpeXdJ3tbEyuip4asxs
HIsbvdEuBrsbgrpxMeE+0XXnC+S/4YpZoVA0IxC0NaOmsecNzal8htHQZ8jYY8Sr8jpFoaXX6lzn
YnF/Ox7rwFh6cxsOy1FdftM8/5DKTMGekOsYxoCgRnlsNVPgPPch3uVTDHh1ERWyjdzj83lKMKDW
BbWOi/ifat6hbEvbjb1vYj56O8CODdwMTNAdxuOIPIhrHS2nEIfMF4MiuMAIOwhZGaNaTvYpZLeA
BjOJsckyIqr/V0nji5Hm6geYt0x3D6izx9wuoP3ujTSb2O4liqF9pIBvCMCYrtIaG4WgwiZKZwWp
h3+bXtfl6qAhzSrySDx14X/KvbTJ2rAgjoWDDvRiAyeE+GEzsA8V3MJ4+l0mZsj80DOgF+k9WBqp
O0SW6wLnGdYQsXIaDyg5mZYMCrTUUqmPZ5k+mZ891rgu9AoCmfVcX/l7cqd6l+5SmZQo7E/po/Mt
gbIP8mhHzpQLsKfHwRqyyoLm0a2TOzf6Ai/U9jBJSnUew577/hLq6og7VmTt0cAHNmo6k7xYWzAi
RmE+Kn8fjlsxS/z8NeL5kVFiS+IHHQn9LpS9JM09N7qMNO28l8cug02RuUWa+qi2U8InQkjkgBgw
F2mFnWQjHLveUPRBeLtlddHoRvGvEkONoQvYpDs8J6+EOall/3R+ub4VC0ijKGL3WLDag8r4+HrL
o3PUNZsngzNTCegmOGXH9P1OXP3HnV/Jh1abUzVeNEiNPownYsfMK+6divp0Tc5HgJZO90rfzztK
Ux36+9yUNKpJcSy5Knppe34o5HzgBd+113Bp9qoDri7gofOuTbYE9PR6zULN2fQ+imrluFIU43Ye
B+LcsBQtI5WmEGzYnx4yhsLsDUltO6KpXEisRQbeAOwr2ibUjOGV2LQ1Vvae800ylX11lX07foLm
P4gz7DzU1p8Qjk7KD/wyjgsa93HPhYbcYV/5SNxRVk895XhGk2X1+1eS2VTeCL8lxBl0I20M5J8p
PZTW8kNMN6Yol6spw170SIIfBCM4+WhRKQ3m2Sv7vKo1CsxTrEPDj9sgEfgdcxgS1eosg9X0khNc
o0pQO0YgjVez7p6W/nSRO1EsrN052h01rkAHiEhiYTYayxg09HFVPvKQ1q5OPA3tj7qo/jbuv0N6
Cmtrp3+BQb9e4aGszccXfKCnrcI+Gz1VgHPFyn5eQjW5C7ASim3XaixvDK40LvCAuXeOrHKPo89z
v/pKr6vhZL6pQYIxPJtkdTl49adVemga7Q155JPgIdK1/oYC5Aaow4z0m52w/ErYCjMUNQ9x4i4R
0bO0WcbfsPQWE+UqQ2lBhwuqtd5zjOOZWAKkcY80xxjVn3idk0ayVubS93T8OkwSv850Gr1mVgBQ
eUGmEJZBv9ZPbnXAGWF1+nlu3esg420oIDgSh4ZbWt8/V7iZeSrsGlmRAsD+WLwAW9T9ZoZ16iHX
bakVbzQIKjSjyBY9k5Qj3Lk8m76Raluz5IvgsYbCL1ORooExpd8i4wBKoU/oPO99Fy2POA3+hv0/
n6l5ajG3cLlGqlLTZ7n23RzoUpbYnFT9KkI0Jl0HUMuyI6VFklwSFqe77+8RMRXO9XuuOPs+9IeQ
I0UnCV1Z2M24AOc4egreiaY9sLx/cFXXJeQLeALDzfkOEL7BCvzlhtulX2ZyEPWO1vklye+w+dhx
4NNWOejllURB3FfqZ7vGS7zOMU0BXSbzd7gj+d8RUNkZKGyXFDMaE77eMAcAArHbomzKaeCeHStX
3nzzQMlwHX+LiKgt6P8BPGt3AYQlfVxiViRB6xActVh2WJrCsEA79Su/dgYgJL+ZtkH1yV9EU3Fk
c1VTJiRioPwxz5FVuck/ECk5hvHocw5mttJCzoGO1S40yHBYcAhCBD1ptiZATyj8i84yRKNePI71
++LZ6ygKtx3fiWYkMu8kRFJilgp9ldCCyOlBiNmfzHFmVaQG2eNmj130M9TXgI+sxuO4aoHW+/hN
rYuLEyLFBLRd908GzJvHa8ILA6sD/NFM42iLAjZJdu/dvIUUVa9nSzcOLzyol/Fh5okUpSnl6Lg6
m2kbufuDr5wCTFji+Sjr4TXisoPYsA5oAkUqGw3Ehk3Zltrjs+kFC6EweLxtBdHU2+K1XXjroLJu
41Zt81JcCoOOACopoBThCUQdVIRs268X/5kXP6WG/iB87RnfzgFsnrZGaxN91GZ6VS3FYp6Ywvu1
CiejiqhEk+eS4x27YI8kViE7YvUh/6RSnuTMOVdOp9jSt2hkbuGn7LhqH7dn9JOOzJVfjD6KWQ2x
MPkgCd+yToFd8gDTImlIJ1bsrd865Kd3iPTYLQsKGIJ1TX+/Z8NVWScdbNsSbxZu+Wvrgta8ChY6
+dfL201n3Cg5nVapz6Tr1KftS/eYRlaqsu+QrdiYFmIrLMZGLRc4sWXj9RA7yVBxVFvA2SEkc6yW
EX3gr5exb16Mb9Oe1qYlp8eKViOZ1xldTdg5+VHIlKT7Z/jkyVl0TYDJssXwYMwI3Tk+r8NYi1nq
YdAN/pFX/TfPj4ambmOTIfWZ012MfCxNQXnaZbfTLBWjt1sn3KtPsEV5k8Ezbrx04Iynji31LQ7a
PvmntpQv5UWWARs3iXB+CtXhPZxKgY8PtAP8Ks4ru43DviI1BQteExf8vZ4RKwAfrFptnpytlpi+
jXS/bSIUSRQ0HcfvBXJ20+1oVygagxJ18BJQKCoAcQuLJH7pz6Lc2OFpizs+BNsq9vRVTwxp+WOj
HYNhEtpm801Fgv5w3OdFltHujHapIF1TEveHJ6O3tdKwtH5NfOxX5wzy7w/i72Dy6umC67rAoHN4
+OqzmKJXbj5z+g886YU70H3V8hgfeiIftOISbslUhajsVAsMg8Fdub38XIJ9IrE67+I24TgVwvgh
/xGFqk+lkUyDFU7WAj1koBLusET9iLsTAzWcXI0nND0jHEW6/x7bC5GUkV4Ua/YNRkDkL5CRIQdj
p/OCID3FBKVU8Ayd/dMb+8pMdTBjOj80CLyRwmv2vn2OiDaByc4agpReWYe5zto97nRjwi5JaVZR
t0e9Xsjrr3towMGeCipZjedx0JDJ1oTo7xJKayHvo92EclV/8Fjpm5vnoppUUQL7F1Hh8u8Xpzbr
A235X5DdqeoCVGiGjq01z+MgsO//UYtnybqIZS91L02YhBYq1KqYpGMGKYtI13Sfgv+AxD0T3+SB
mlH21nUlYdCBWOPbOl22Rl7VSyrxSgTGRucJHJ62nI7l439LqQc/+10Rx1VjgD/A7e2w5e/TB0Go
P9NrZARY+LrCKD4nx/6YGi8cEwu3WK7Erb3cLehuFlGDETUjAf2kPdE4Z5/w6qacjHaSoN8U0F8M
s/gkewUoiuhocv0MowooNgmn82MzUJrEXgI3wH1O6gVXuwonUZjP4bZe06iGX+cub7/fVzfsmh+D
CcrX36D7AvcQyl2HNTiBigKqorBVcL1FZIC9TUOVQKJaFNl5tZnM2qqRyqNfnJutjbc14A2itKq+
OXdKe5C0hh/1ryeJXdp6NkD6fy0bAr0xzJKcrnUtp5JX0E1WV1h4eElK83Xro+ds3r81k7Hivx8z
W3zy6A2VaUmo9YoM1Y50N2pileTlH/VGv1CG7VtwOl+cX051hXKfomyw7zbuRdwtTBm/dJhfsh3w
Wbz05J8NpMnYDoVo+nQtnO77oEzUHgyqAbZfr8BbLRkOHVza0H1/Mi+TKk1Wvj8s3VZDu+7lniVa
0vuP+tXkVsIajQHf2hcN2AwN9RTVbvcNRx5sPQLBYt5f4XVBuvJd9e1+y3jNVz6US6Pm4hrBvTxp
tEQlknkPaDiY+nJ+7kbUx0PnPE5wVNW7WONoVp1qqlpoi1wMqMj3UwgapYOIWUadqEj3uwRARdcd
7nucyO6jC6VzsANPF5ToAut8Q/5kX+dY5bkbD2M3xx/QVCibDV3FILihojuOOxzn6KFOUM+uoQc9
fF10NQwqP/cm6u3UtrukVXOGVRnO6PyjyNJRECM1QyFEPz/RKY9E4PsQ0RTS5dUHupEWxp/45Ods
m6cW6pLwS2/df/eNnFqRRO6FRC1mml1udkegYbuqvJnleIEcbudpXarDk+9W2BIUVsj2hoWUygtM
FAZdLSsNX8/za6BUK620gvtM8VwnA757z4PkuzkqZZ2hIRKyg5o8rsbkpZ0FS9SCbnjkU9bwTeJQ
Xpd7bdFO0l/72bkxWkA5fUZaL3xaLkVaraidKHAoULSR6ueWs4HwSL0UJDVuZ+TU5l4+i8uVYNdp
E0sBPmOlxai9CvEpxbB+0szgz6VdI6f0jCepkEws9HwtzWxUh2acd1fmo4jyXfgpePDW7f3gwnNx
g2vggiWlumcxipmH6u3VCIemCJNgAFxYVcTQttUHN1xBOzeXRydIhHBiI1ydZD6CPAEDgsWicHFi
D/JUl1exfetRQWXtmDWpXlD0TpnJ5PZv5AzHaXvrTQQyClQ64w7cXYuMeLqPXc4AVjgTWlGcbCAc
rTtiBonAZ+atOLU6eyzJgCm/dL3JZs8/8snrZ9nxofltbqzz3XLE4GALJzHNib+Jps0+myrENccP
fhJ0dGJNVT1H31cXQJSddstYvd5L5QUvletCEvSobfDZmgbK/Ue1kuYMSEWjgx2QMlBmz5SydlPS
LYaEfdtIHQKcbCZBbuhK4Xv3G5sEvrao0h3IZEayfWawJBr8jpawjKvzBq2+tZ8ZzvkJR1yhwnt7
oCELxPJcN5jBAqXCKy6Rlakc1M7riCDyt2ZJClmoYHWvgBy4MBeh8XSFxGMfneNdDqyHEQuiffu6
41YG15PGBh5FyKWJ6u75BuRQsyUv1W9vsbGivViHQbtKZQjoCWKYht0/rFEl0SZnJNUSMDedSyvf
XV2cqm/JKolT7GOP7T5FDry1ynlS+X/pqE+3wrk/yyF4aB3YAtP/Ffhd9/6jlEkbIhGlQ+z5jQTI
YBPEeB8x2EINMlrr8l7aZsh/gN7GYBTQdgCBIG/XZ4NLMSyfs/6kviVwcVJ40oWyv5Oj6/02fvmp
QLmLHLjIrdHXXUMzJ/wpZIbhXaA/U1haY98UyXpa4a04UMtd2IZIQo3GS+9YOAgpno6nCw3eUHfT
de00PrrIBYRCO5HkrUp++kZB4OJm3XaVM7pn7h66jk47ImaKrMhZ9122bZUqBWYF3laMUB2iMhKp
Uz0ZYbcV7y9fsfQ26E4X821vRHLSuxTSbGhlkA19C1cVYbnug9INYds6qyzlyerGUTkswJdHkvfi
vK25wFiUYjE0J5tCboGVIKNdxtrHp3tf7KWJndub/NUXtQiwJIVgFvmBy6lg94Q+FCgtmoMpLQu9
iYQOmv/bEwukFNOSk38jrUAfsWzO54Z3ZSiof6aY3e/2ES8z3tGFcTjb39/TJgrvAjUewhZlJxWp
IP7au0qx20BXzi8Ab70HUh1rtNu3yq/2PgA5ZXWrO4w/cHDNJk3rAx7ApD+lK2YszSRrxzmKegg3
EmZLHouG3djM6uyzqdKzQG0k5AjVEYfFtdW8Z6HwUIwxFK9SDH0xiBXL6WSu5cya5wA7op5RdA+8
oQLiM3WutW1o3N8hGK+5Waffu+ZrjSwA98RU32dEVCDQ9tCAbs9ZsyviBR0w5b5oQ4kaBeOihFKY
7zJHQoMX4UimM4GsjGVRpMxZgh1+sZvEW8AEdHW0hbBwc6suWBBQBVg5NcDE7enbEGnI5vZyzqE9
FUMdQmOklNl1CTTi3d2W45vOozbud38C8VRxdQx3A7l5B6ST6kWgbBi+l70+fWF+M9Cyhi1aKJQK
xC4TPtisxLeq84mR5QlebRjlNvc4ZkoTjsluuvk6BW4Z4I/YYW0ts+ZonJKhW9ba2MuLJozdYIzZ
CoQ0myDanQh3RMu97suWjKzIyTkpMhq3W1WyqIANNQAkeaj9WwQuO2Npg/+b0MxMRCCwL8jWKntl
8fxpB/vMbnsfWVCdeHA68qLp7KdxY1r/CowGDM+CiJiBG0rBvB4QpFuyBEta5x7QNk1i3gQK2W5V
hGtb3Nxe6hVHSv2jcRL3kEr+3Rq8nCPNw267tt+qnx1dT96x/li+ipvIeW7eos4WvJSiAw1eW38x
YtMpb+jqGVzAZtZz77mBI8b6Sjh0XSdHNzLElp/bh8gmtFTnOR2TkNlNKHESxoHhZqLb6/WEV8pZ
m83rPguSJE3TA49MrnGIGDMKEF4c+zCe8OoeG3NZOyZnie3BBZFy2kSI8iU4ddaAg+aL3oZ89m7P
491+6ik87b149EzDz1tmvI7Gae2DGufTs0vYCCO/sVBluCNGkH9xOihD177ZvDAL5KvApSTn8kdH
Am7cwlFwcX2IMPJuPfRm9YJ+ArsW0rJ92bw2c3gHQbP749OeoaUc5GZpwRtjU110F5x9RU8oipTj
KZ5kxpvzFAte4fT3fDojo1zRw+n2+/QN3w5VDMR73279znMekX38FCF0VnHunip0cS610UZ9g0n5
io2aJH96ELqef8cpjm+MStxfTCEY2lh0f1FXHmZAcyBQPTCOByvx2bB0DeVhkM0lbLaLiF+KqCBH
J0MtnFJSfr+HjNOUKOxoqaOR5PwhizI8I2gHCq8IlSOfVw9ORzdCr/Y+4UAWEpDTEQeRdfGTNVWp
XU77HvP1/f7EtpsDQHkMRpyEevttOp5v83M5Ikdaxk1QP0A4R2jhSh2dUzUG/lD7vzr9BTWpIjYm
KMl3PQgmgwYpS/5UW3A8GVMNZxnUtUZ7meuVbhA8TOylGfuP1TLfMcQraqQXKlgvEJy6GMIkLxaR
I93C/8Ooe/uNVUW9VifvuyN5U0lLSx0Z38EMZ26vMF2AtS8opMNRxQ4E7Gib5nLYNgnIh9I7iDJb
BbAwXasU1cnqFUqkOR+gSwi4lhjz66C2ollB7lSsYSqCHIIFPvDBfIypL6S5jD5oV0xKTTbIFms/
yGgrQ7jjBSlmUtoUIisUJM7LOgnXLGkLdIx/ec6/uXtafrznY3Iithb7tZGzIc/LHxN4O/W+/h15
2FBTdHRzrM0RRidHZbhgQj9wmDgav25GfiqntMEr+9IHsZCQ3aI0NuIMDmTVk6DICcqdy3vjNtR+
1xW49pBDjacHVBvIsRnFioG+HWB7vLkJjAlW6m+TLUOSEE1E+9HkqF+y+YPZDMa6uMhRNEUKPTIO
Ba/+8j4pRy5b02Nd89SOMoqHuDa++QyeeIKYctFz9lYQfIete/FCyIim7m43BP+2i5pUYW/CbaYj
31t0n5zhl25hIGd3IAr3ifda0i5wiPea4g5lkuRYQALA1ktaz3/wAcx5c3QQuQWBbPyMH5hCr5ma
4t111Yzu2NEKdYQfiBLj9ea5NclhEboHlf91YMxsE+e/C7tZ1o9+Lx7iLUmrx1yz0J6DHWTzd4oD
T3Vaoy5qETtKCSdfX/sw6MmjnJi5DDPKdqUCHC863KVOEsPtOIrLWe3/C3PVn7X+kNuDh8UdLae7
kimOK4lr01ehCftyAjsfEpCc8uK5nyGhpmio0Kb3/vDX4tlx7UpyzEHekJ3NCmrww17XRohloK2n
dLzeRhEaIUCHBzAmRvVbMNs8RXVQMlb5s8LE6deDY+iE9ssecEM5y8pS57MW15zywfD60J0Zb8qA
VoBlzuqGqQzusyczbMJfIYQ9BitawvhUrX44/0DdqWPsZQNcF2sZwaEULKLf5jIAP+o6bmS6awB0
wJGCZgSWQi+3vma26NOUUtf3IB5wIkQ8V1DLGSEe8YmdmkBXBxUGGvZNJpsiq5ku5Kks41sKGkod
pJYJYHXT6ARThIULmcW1Aog3UBf0sV+VmLV3NIWKF1mOMJOSFc5jlZ62Xx1N/8UwkPU8gyMULaMr
jf1yHBbgDtNXvQvaesmHhLAt0hCpHVi8Xhv6cEbn/UkUbKyFeF5Mismb0QYFO0fKDvE5vPtJWyr3
IsAI35Q61nDoKgUEEjRpnx9XEaT+IKOgyRwgCEX1opdaKcNzAysaIjPw/Af6yYZvr7THtklhEHll
rNjb/bgd/ummVvawydirLV4u0ZpP8rJUnH7qqX5LUN9hMLl7L3qg7o8487Xyt026SKMsemykuOSR
f+e6xBGMcdiAgkmC/UWSInYJTZ0JXKBBu4KTCCQrO9NlPdnJK8dfJugG1QKy293pDcvFc2H4sxuE
bBvwkbJy9ht8bHuJZLGBJcMxHT36wLM3x3+bmrt6oS0v4HsAdw0B5AXGLWbNhDUlNPE7ZkBUryXE
1YYwaFkgTNfqWmcTYswLntbuQCeKXgsnxk98y2EWbnmKzO/7tXe5ysAJkpqv1GiHwzpWam4J12WH
AVvOyp8eAZRJBOO7PlErCkYQ44fQShEkblj5d2It1GKZ4C5BIB9tyfh5unaZB4vhPpZtcj000T/b
yyWfM32TzQ7qzJQxhs3ldrw6aRezl3XPfWX/+/hhLJXoRWR06jgPTaticCFOLLdZRpNATV+/Njif
zqJKdDgCr1p21d73Io3D4FP4jdixK39G7/0QwrIJN2NM8Fs1eeV1krz76uE13a82n3TJeWycjQMH
5pGyX1XLrqK2vwekZf0W/qrmCGkooUvkbvaTIOYv4NxQNqgBGA7zCnixk3RXLDMEfYIfj8PdmnUU
TfgH3irDwWMdb3ETrJiED82x6cyLsALpcZUimDKolX6SOYiLz9Wl5JmGPj+N8+1yuBruTWnZ8Bl9
Rez1M83xsVQheTkdO1cZHncEtn8AieXTXgO3QLHEbeep9ZvAWukJMSPZJBMB9WGFvlws0fWooHJt
gR/V3iBc0y0THqrCLiw7WfNXbYJgHpETm8mTKkjEnY34ukBlUYG+IaYvXxgNb4WdIqifPgTClvOs
/7REyhtX2CIblVQpTiHFb9A86MP6A4v5wgWxEwEk6RyAfIoYpeyl0OLIvpj02MQkxNNTOD9F/yLc
dQx3p6k0kScV7Hxbt2Gn7Unc6b9XBOqtdVEbVKW/1Nqw78YLhBq2hpHQAtEuUtH6UuBsmpgFud27
A+52DtuZ9lGD23JwGqm+4Rr/hd90e4YBJKDxusXnu2PDcdbRzYk/mnq8Jw0bhGB4UAgGzhnwaBch
hJPwVk95Zu+ev49EJV520Z//zs3oDlpX3vXcKDYkvM/GbvbQyfmlvDXJTO4+l75UwJRWluesnr+B
Y+DoqSs0aaB/cefSH/QWRjDoo2kTG/rypwgs5t/gldBhF6gLb3vInRyoSL15iJAlI7i9PXdva4PT
DWwTBFzBdPlA1uhatGoej64MLwPXvqrnE8HkTuWay79OSl+A3woA/KnOvkFAS1wYQh0jXXjQdEgD
fhasajN8p46D7076Jj6BAaMpn+I+wOSr9O7etOyURanc42zdE+56YlBgYnIAcLb9nsWWm6XnkS3n
NLbRcDb/y5TpetnPxvfQ/IgVeldBICGnO+zj8+M/u/UnodMV08pyV3NXQJaGtkJGnzsEv4XEGlE4
4x0boTutFw8F5B5NxMc4Fg0KPhBLfiDifhsAj9PF33VFd3yp5jEy+RBvULP8ZSFlkXA1CUlldTdg
AzazgHWwFcHU6EgZFmSjZcmAwy2QaC1mdINXsP04y2sPS9D4fqaVNvnV7macDYe04+z1q8pwdkIb
8dEjNr+6U4t/a7hijTz8qWcwQ3mQjcGIQePn/nkFprNNcRgoXwefZEAtAdenQzRcZaxLjdGRG4AX
BEA5ZMVk5nm2mAa8q8M5nf9HV0FvjWxucre5M8QQ4k3GBsEAitL75KO8XdrQPZUH7cRI6x7P2rJa
Ei5KVIS3B5hr+WabvT3F2/KpV1s0ZDJ7yujg5rVkjvEwAUV6UmXB+XvL+zUS6HZljSPfM4LVfKKp
bovD5bruMXxgG+DCfdOjKKDyxCTRnxnzYNcgkoC2xgcUQKYPa4aqw6rgV6ytpY2d1Vjf6mS3hCJG
hSGwWE78z/a61iaJZIhfvuI2uOxw0nypPZuq5mpO7ip/duwWJM/4JBTjbb7GE8Dnd7OFi3TtV4aC
MSArIAJzm1jtqQpyBFf99z0w/a+a3sOnn7UtHjrx1RM21P0ZgHQ4TTFr6YlsMBM7ySYMLMz/mr2O
QLB9KBBYOMHT6ZWMqzYH22hFkMdVUawdDLapYcJ0mo/gnWig2GcN1UpzakJsWatMOI1hZJvBX6mo
sv+WKQ+Az2BdLV6fkFEOCw+Hl6VJ70pmWA86YRwBZiTCxrbVElEqRvr+ohX20KjmpCwbu30vydIf
GYJvgFlyYZrOff53xX993YVPVPwf+AYuRL/mU8rAA+1YyuitiCsGIEqSzcMlxOVJtWZKARQ6RiFL
RFDLix7Kp8k7XhuNFCRxzRHrqqCBN9cAVmBrNiVggDz0KV5EGR59v68QUqAiDD7Qb8q0uUDdaia+
7wDxAZYd5+sHICGPFCNg8Wo9rYaUIGeyMOAeKUIqvR6qMw7DezD5aI5xcY+QhlYDGBVt7Yu5JPJf
xMKfAGvL7fVLzuX7v6e3/8F4gn3gGu7xRl3B9f0BsxUa8WP0bToJxL5aR7akzMxGHDIYeSgy/imD
X+QhkEQVAUnuzTbt9RE5CkJUb/rNBWqK17bwqX0F7AtXsgM+HQoiVTOtCNaRB2N0caiyMPFBmcqA
arwOeZmk0gfh0gtLqu+aYF4Gbwoub9qE3hG3bRGJQAzuV03E85FljoJf6BwwRb8YHJfm+7yBifNP
LxUeh9xxhrdbPo5KRfOCx4yXnnofhQD5aBSEbRe0J2Q3BE409UP08dFCG+S+tm4FUZoF9NEU+Seu
zzlweg4Q5keJpYfpnoiDSsrxrCYIavnhngPKeu2c6TZxhW2Nwa0TVQIYagHDRQJWdsIbEq+/+An/
/N8Bt1I5FVGxXMvp8wAbBzVWKqiwKYrCHdfYB/fmtJ0zXQVKac/aYLwWmN6NP9Z+PO7+MM5FFuSA
sg+J5k2iiy4diBm5WYvEdPkgosQRNYkJv+u61rSt3iQbytG5+SnGG6Ou+BC42YUb0Gv01ixYMQMS
o7jMn8oQmuE+/cg+QtBRXdSblM5r/IlxmpelxgZaMqCmE9qZDze5+Ff3kWoGjqrU+a3inP/Mm13z
AQnHbCe5mE5OGRbW2yM574Yhv36+3UZARYVTnMBSeEd3PPAkCBsMPx2Xk/5uFl4/uU6nHx6wNYw9
4Qdhs8thWLv5DA64zyX+Zr/IVBNbtHNXqqzAJyqlzp2ohP+o9HnMG1Kzu57CvQlD4qfhXZMCENU2
wO7iggaxDifHdNviKjniRtIVhnOmEbh9t22GC0bYODlgaJMXEpr6+vaw0a6o3MMYxFke8LC3wDdL
Ph2jT7Vxk77bAgCmaQcKcfyeN/b58Yta9pZMULtDI1gVZNazuEvfIt20gAlK2rvIW4JfYE3xvsN2
96+PgWHFQNBCHbYjHnOMtU4cbk4VhEUm6PMLnOYBFjF2aufyEFqpeoNjNmPD+VuxtZkAJglf8b0h
3wwDblhIBm5y8YUZoqK0wsuC/XzoONo9qfmREaiQ85ZPTwcSN25ZnbG56NQeNPUOkuTOHNLydZ8Y
iGBnwsv5V8qWq+9U+DFpZkKPKbKjHESqysRpI4P4IE5v7gXl6wrYSr1uLEHkAmEMIj+WuOccAc2y
TBfqQyGoPzZj+TzD8YFoPq4C+sAJ5LaNU0eswwGAb1mrWSGGmOT5Xw8uwfGL2kJnF1eTu362hebk
7D2fBG6BkzhixTevQsSJAUvyaSwj4I6evLTI6kVgR6cgRAvrP1jmk3X9WO56SQ53VLotaSF13hXv
H5lTomE/Buu4FQvWNGPZuToecUxanqgG4plKLMMfVQ7DKQKAouNdual3qvPPFYXq6RAjE6+koGY5
8frCHS4bqX8PVO5De7vuxpZjxd2Kiness1Cel6E+mDu58GW43BT0enjAgqiVTf5qj34n8KhOsieK
B0zQrCbxF20fCGcok5f3bwRuPdgIkVumEwxWhQgPPYlHGDxeLDRf0Pm3XApNOKqQzOudiQq7e450
qmX03TPvpoNFzp398uMuAraSJJJPpCdDyziNI5qsOo5wZf3Xz4/oJBgW2ugbIE+Q8RwhzHwLIEcl
+lAkkungPImlYdd8Zp90WXMwmmnKxY5DjHQdhA3yIVEvsQiaP4R4N9SycGe/QqCvz7V0Hkqt6M61
PlCses1VQ0op1rwBtxr1Fk69ADg/V/z/Qvam/8bxUWjp2CTbGfr3Mqx2WgZ0Tu55kGeI5jRIRDLp
mpJfqHL+KWjc6XTVWikaAWQL2QOXu21JuUlhV71bv5PSs58iluwujEOsGt9+zATgqwYWq4rfufRm
9+777431sRVD3lY72q4O79/c5429zea4JRIVY8ptQ456c0mFDp8y3f/0CxOZhRKo7JnFHqLwMVyk
nCYSec4Ge+rmwoULGVuB904gYHO/vzBl7MhO8bMVIzvV4lpBv/Y8pp3v2LNgPrW6QnfY8L80KIig
AYeXFTYxe0hY5nLqxpafSMYbNN56Hgi9IWS2GfzYATe8v2o/rccUAmqKM8Oc+CtV4h/Hb1ZiILDT
Junt0uauR9tq9h7H+HxqvAIskphbUbu8dYgoO9jXvwss4eS0zuGk9ikW1JsK/qNAKbBXz7+32fDd
l4PJbK9uaKUv4BW//4l/L8sIaoU6lbm7BYR5Il4DB74ej4gP+ce9k+GRzgdelYR2QRiY6Xp7jcP5
moEmmASSr2k8UTbvFaAvf5+95GmTBiB21jtlf2OlEgatc6nfBzNhNyZC6yXuHxuV9NKZ5XetYOi9
xR2YGSRxuISOavAdjqrK8xqyXCNDOEdPo13+72KPMzfZleyv5tKO7nYvfGcSsXLDyprOegRx5evo
Hy3x75Dpr99ZlOPJOiR7IEfYz/uIAfnTaB4uO9tEB2FhobcMm2VXn5E6c4yvSBa30BpsquaMuFFn
XAy8S3Swyq7uQgm3ehFrOB3UFZWIewiSO+vzo2dNMxaGtxSpSit8XM0jHiMLaITkXxR4Gnazv7UH
ESktmAhyjRXDOTCIREn3jeXgDgZq7MIJ8Ht3Blj+YuMNA3twMd37Z8He5He01k47u80CycaeoteQ
ZrlI+c5RrBfWkKdxj0q9CIQto/Pluy1LRQitk6kykkLZoZiM+WT/7TnpauYgJy3WXEtdhK80d1YC
m5M45uvdth53z3mQrhlk2YA62uZEnPgwC/xVACREgk3BrJWocB6x8GishvxAZr4S1ZSyJf8kZH0C
dxl2SeLj1PGZUhXjiZkxwVoq/JGBR+et4hPr3i6KWL13FEtokWu5kHpjZWhL/8X46eO+0pAAC/jb
bP3QTeTbfMblq+YhRELsADd4cCTyIS5MC21sGhwc5A0B4C5FwNnXffZF6C6axbgQSwqdNsBCUql/
TciVH4mGLxOPIgnpraxHQbjxr9ABlDVUOP8RSjPX+CtiHve1n3VlHwmGlCCWP6ZiAONLpo/zG1zo
do2YvE8sZEqN5nOAcu5Rokm6Mwz5HPKX5rza3YXejxx2ICos+p1vjAU+JZGzSCU941bOb46X5l41
IPo67xsxwc/t+7dIAPYMRBTZifflaxI9DupYpKRn8ICxsyywXAwmnISMpBvzg7lULxfx0Uz9UXq4
pkHSReO9lc6iPw1gmxBcUz0PvQoYRsxtSfq0FXpD2BtOHm1UxTArjqNX+5sb5ngtiUVQoXQrEvHZ
j9HBhm9b74eu9RhGMEisoUuJdtWmdvHNIygVPSRlQcPxf/6nvOZAC9r7KT2KwLG8iSBegWzeavIC
bGciKSW27WHELi0npxeltOVwvyrP3+Zx1w56dj4ozftcF6Aaxas23xMJujAC3l+G1xGZLYuAKucR
im2sVh/ehDPIGqJiHO6qRwCk8gUYoWA5L5St5ZGHUXzPHbGl9fCehKyWr3MJwTl5bgqh6qO5M584
wOfs2rR0l01Oh86CHJ9+40CQWywsKIxB9MFmAvuxbLdUpgxHyS7hN0Uim2yNFOm8OFqXrCduBXn6
pqVtsF2PN703OWaeSeDA/RsySSNUrUa5ko68jWG49YNLLGyq7W18dO4gefhJR5Gs0o67OFE5dgu+
W2kUvdKyvvv6mvzmZMzxB3xoTsyWdZjLVYn2dttjXa5nBPd0R6j+E7JyPQtq2b0Soow1AhCRC2qj
jk1mvnFxgAJwEqYskdqo/Zue6Vb2uLEj49j0Jgjcgr2nY6zqb9BzQVDxIHGf4azYyiO4cPQhZQ+J
xwxjBkI82TtpXywcjzhWdz1Y/AOFcN+82TMpPPVzHTffzkOcfObzW4QHcKHYa+ZMsD7Zd6S4He76
KQw/KWe5xxT1LXv4DuUaxiwIYTwSOVSdjdoYiClq/JO9ta9u6GYrYyqudXBa/zTQMUge5BppTDb4
1dgrFMW1qOk3Tw6on2pPczMzMoxaGhnhRu/CdL05B/IjQHKLdnOSXQSeyNBxKfwPy7qldUQeG37s
gK0t3/S0tfI7OElOvROi4QDdhz2avmcNG9/lP6eXfWmgoLBoTnn2JtBMALSNbHfQnwnUg7fxA02q
88TSs08X1v1NSgbwYrQ6dE70PJD5RqDwPtbLZAAfIlL/q6QXBsKYPYhyZdR++LNieYNkgMdzVQ/m
J3lE9F4Cl2eRlRmKbq5eG0QJH82GwYZXXbLt2L6wwIOSvD/V65SxgdhOgq1BdEBmIjYdTn/H9qJo
Z/oqTh3HpJjenqYLfN5YhIWvQtKlzBiFUqWfNiWVs+zzbIGcsf706ql9aDTM7tDSrvEWfKY6BEuo
LC9Hb22tET/PQxl5r72gxpYTK7GDcO1jBYx/j11zMDmafpVq3okPe260Cm8goo28fG7dK/zFKzdW
6FhC2Ek4WAIxtQ6/ZHR/DguHq/N7ptpq+ZAXO+jhujRv5KJWm+xcabyS4QnZLcJs6R/Pobp4fIbl
eoni0hV8FZ9w5phh7IpEiAB4cKu9bJefN9WMhwR7qEaOvfGjK6GndE2eoywmHw2iwAKpmbO1bH+f
4aeZYLVI9Isz4yvIVtPEgen60tfUhE6ttlWKUKOgoah4dqj/ZvkDNtDN5ohcOv6AcTA5s2q9bkyP
+nOWFtYaRTeiOcgSNVlV0GZco6qE385RdSWUb5GscuoaCiQtLKotp3ebTfRZgyGqCCDQMmrYqs+3
jQ64e1+o5jEzlTIUAAFQoPDvsN6IkHCBlaqCWr0Xb2BU2B0iXndXU9xttRDz3DDJZOzZGaEaeK0D
0WFCee0Snn3JnPOwIIRYbQxgqmDFYMy/sPmOw/D++ZzghLknods3/OIoHocrTwxyRv2ebkW++uyl
SLciOhQvcHLKs5QTSNSt59L3CuNwjfR0K6//Kf0QnBilayGzHfe6f0PpXKJpmefi/kUIhf0IQGF8
p9y6wiqsF9RfbXnvBfCU2GMD9dBB3jYUauo4dre8dtHOsdGfoi0vrICvBfCMdUvi+dz75kySJOOS
eIbqnet1js3B6xrlLGiutJ5Qlr1ZKx1GpOgIUJOG3Ja60rlyzYf/ywyyF0HYG88jSz9NBZUXy6pE
hDoElzqzgTlVOvyNVCyHeFIXcKdbxXZi2mvPQrrYYlo1YhProioJJz+AyJs15EXkD8mt+HMJch5c
LhW+BZiwY3/DFhSSCIR2Ejpvot0VNGgxxwa8U1DEU06q4ypuSom4v9Ys5yOTda5XyPXGkMXakAr8
jIrJSQwdcyFRoQ5HGyFDS9zeBhcdlIesXq4uERr4hawNPzNcQrsfpZ0RSm2EepknxXqFTeOruENt
oKUdMWN0HoJSmN1R55hwEACYSvoSH+xMiF4NZ9K8Eq4ymeA92aZBUIx38jSO7Oonx/qbXFpKiwjb
HRQEIS/D6s7yiCatShd5HcLDPOy/FdTKlMEudzBhsWl+Bo3wYT7DKJEERMLb4qyWIfnR0uCFsHQP
+XN2yaux2mtejvuZW1Mi3JTurij/k+kydi5nFE53x1y6HSpyR4m26rZtB1N7zSeJyJR3WVCMrstU
ETwNMRO3lWPouYbz1sualplQtsNVdxhb24K7aUKvqbmF6LMa+5Ur3FPK+XN9BC7DJ6420xdGGoRW
dEEDvrd2tpInypCAlMr89fb04GKm2pYerkF7FS27C6JzcrD4FNHHM2i7SaAJslD+2Bn+ceEzIW37
nOJlDbb0W5BhRKAmA40mzSC7hv6TfY09oERedwAD4p+i30plL9gn8QL0rY3I/OyG60AWeTNYvYt7
4bDDcF05D89u8cPAtjfQcXwD5s/89sNdJMpqG5dwrhgBWpzdMFm8ncC3vmUTtSED7+JW8z+Jbv2q
ckag3h4zLzXWBRtraWx/u48yBSjYQOrdEmhdkLd/a535HJ+fRwi+6+VJ4L2sywB2VNwekU4xzogc
Vy6pd9kFQRlz8DaBvBG2MbjfFHYVTxdCNXnETrAYa6dcMzo43Er70ZOuuMlRJz0bK3sawGxKSJK1
fY6eXF/kfzsT6TfM2JYmJAoncQEO8gfOU8XUzXGlo6wDiWsTG1TiA8Rc5TIArHFS3519Ir12Z4mk
nrmRgy9Z0qXKHtOzeuXQyVOGXb48mWoryDXm6W3tVZ6GkBKqCFx5Os9Gyn48Dgl4hq00HGmmT14+
uIjbukbkGSbdkeaHGv0lDd+XtaCCTdG1aBVX7T4isdNRxip55xMrzxyWLO9fnJky5HOiEM8YsJKr
f7AsTUo9Q/99B5Q8f3vQ+a5AV9Im9KRC19RDQDUQfBCLdfxdKNmYKqxpnsMd2bgNqIKldaqbKimC
ftHQXNWwp1Jdr3nr9oe1NqwRt09taYa00RRnD7nNep7LkmzkiOwktmj/9K9WGUWitlA6h1QlWPUM
wxqPfdCCm2Ubh3S/fWfFfEKS3gSJ0SvjJUkC1Ls5e8y5fkPSW5ozfIk27QK+uvKi4ltCzW2yuE8F
Jf0LmZ2sAuh97UgW4cJLFZHKN1zBfIT0fnX3ZpnCm6fbI7I93HqF56+hXvT92O30ZR7O1/6sQmts
rR4KhzrbU63xsuhcyXAYP8tDPG/fdScy/zd0lhuYV1+dW0cHCp39AsjoeSJZEIQlXu3J7OVKcOuX
vRAXxrbNP3TvlGZl2JEnRsU823jBBCbWd1854Pok0Hb8wwRt53Y7QNdHrOjfXTor95nG+ZVNRJVe
HGFUmo54vVZhcgOSljbnI+PCPq+EB1vG701u5wJvhOCn1Ao2SbkBO+ZvmeamW33P4tD4mWoR53l+
Zqrap0bJ0NjrHKE6ODQEJg8+oAmrJ8n9KEamj96hb03gfT+VOluBQGJOS4+WPlmkYx42Hme5x/yj
uGIktVW3VpG8hAhCqPhB0abd/AvWhxF5xB2iHhhmvAAHRQRdtBxrhPJKUpiJN0opBhc9nimBWbur
pX6ZwoRcFF/4Nx1J9kew3wb40ahPttuEPOq4kIDVfP1EXW79xHgWgWpCQEGiJ19mlr6n6op1EJ1e
vGC5MymN7zGtimQDtwX41gZfN8P2h9bCW62wUAYsRLSoeZxsN5GksDgVkiAJZ2frktiLKX5mc3/3
N9k5R/z3zNfX/fUgiSBqaZ0G+cUkSaBrpaz1I9gme+F110CtL8TJLxD1UDiwAYilVnYOSuAi2QEh
vsLF0WPTIvQhLufaQBgYi19mvlWdXugyZ7OHnFAeeCMCnLIGxrcH2Z7lqTxaV/GoJTIh3NvoFFdB
eY/ctqnJsanviCn200XYooC/jfwrRZ8se4dFZK5djSyEF5yM7VTdOQ+LFThivVxK3a5WH6bDWzX8
GefH5r6kX067u0xdDXD4ZVJjyDfgcP0eLpJGe1l2Ijwedm87iJsOktKNfbPO7EVeMS1Jw1jQRzoZ
feNYfrcL7S4SNC3pxNcoSv035vAMF2L5RWox61MK3rtvx0917Ydc0eN7gHI6uHTCl+C2FbmKEXcV
jMZ6wWRId+mfo3Rk7FM0aFMh9jVQFZMdl/4bmzHXeCAQWIWnpbFujEIuVcEeo/gJ3MqKoOa0hD8V
Oi1/slhD9UivtsJnGTM3/heORH3aE4WrEY4uhLxS5uaidEO6kyI2ZS44DbPSXqSBtsJZL+K8cCa9
IrvWQuCueGESzovpZ3ikIOv0ecFM+FJt4k29RkMEnU2v0LdNCnlYRn9prIxtUpTz8U7DuJ5Kuq++
3rHAXQnCyzP2vweg3tJ0ELnFUFBREwcGjaTBclS+aJcZE7Y40PSSY/++Rmlzf7ocB7ETaJ6Ualzh
IDWWvnlRxmKQAG4OS6xrMKHKRukx/rI2kYo/znbbCynQluCFzRvV90HV7GUmNdh0aPw+FFPH9xLw
cSLxQtRTQs3+5h5EiY1DfkNNZ34Nafgqssk7nXn/cG0c/lxk+h/giaMYH2lfyHvOdL2HS8/u6koS
jjOLDZ20vODuluYgs65SNUgX17BHfUYV2Iu+/homg03bo4sPrLDDQk/J8Db3oPk48l5Mk2i+ZaIH
YIz4RRmWd597/LScgX++TqwKQdVIdoLvuLiQ8xXhDqKxS8fs+d6ylvukxFAo+zlClZi0v6p2k8qV
mGoSSyJx8lyTsDcI8wIv96HJl4JT/eAP2sfpZ5Cw89gyOUApoX5fplx+1zFh1HXuuzJ3J6RahQ86
55clx++daWoKCoiGGb4JEp5+0pmb4Hm1L+BE0pKCEp5l3Xo6284d1T22K+W08N3ntWL6u6vwvP1l
6Z3OjI6sPaH1KAuex43lpkYB0BSpX9yJ6uEESpFb63hvCxEuK5AoyxSEDC1Fqhzb+2JJxkKL1FA+
TP24vK9l37PtQMHLPGTXiiT+1XWKeq72wLyT8qITtQnbL/hw+PS/VnBh5O5nspxzCtDZbT35cMF0
p8SLtME0Mv3Qzryjjy2Jh6k0tveimLOfRf8647nkk8ESaXLkqoBHxVoApmY/ftEcImxDQT6GhfXN
VRftPh337Si7k0odL5dIvL4pwQJ8EWEFFzZtZitVz6WLu59h4B9qJQhjDIm/g5izEbk/+PqomUkM
sBXTzB8mQJ2jvv2itYx4gEthSHtsGuF6OwEC2lPr3bmUfALO7/fR2iiIDxcn174i3nSGIRMDkUtk
mT0B58BQaI+Ls750g9gzJGui6fHAB28whm8w31b10VYAZNmCDiYY18VPyw26soF3XD3kgqykDXv6
QQVRq3aiyRh4QQ+u8asDYZ2Qf42L/4GfqzEU/dmNry7Sjx1fx1WXZEK02DIXG5ney/I7GiqSuEc2
hA2jPETKOaokuDKndmyukk2qZrs8sM0cyLpUCV3nAtbvAj0Ttr161ignJGvqB5AxPhpP+jBWE/jW
9YVuCdp4Xc0sY7ossKoSNPs0kLQE5YDwvV/hpB1xFZX4GeF3AtDQ4JCuPlEzbkbDN/ufeX6dJK61
rucrFGZ9lCmV+HHNeDm4bPe6k/AIPgEJmq/eCyAM1aW71F94/v5R8z6wFgBZUI9fLQcoMHwv7IT1
D7mceVCaqlvIzpFHtbOAeD4/901NId8GYnKye0q+ztxSPaTRv/JfHknd348cOW6QlK0Ze3o9qYLN
4pgkxajyfniPOgblwyZYf16IkY+nvgqGB9d/Ab6waf+KQ7n2eGzLKD8IcXD7zdexJYwL/MQZtHQi
yzk71nk8SBj2aSZEhJ5z9ePhYkCGDYWYNEKX1JMv2Jn2xA7Eo8c49btV6LoLC+K+pkfe7FqNM16X
rJ8MLRImBZJA5mEfSkU5jLaj+lnHcSKkVzi5nXF8Zadw0c4+e1y3pDn66/EwG6qWkwY/ZrV54ri7
TA0H3+0BxTk6tqIXypmQEWczjnGvo6qgCG2ohjkYqrw6SjfEjsEnZ81NcLXkyM2USUGTLFm80+7o
ZaP1V6RrC/yOXKjnkjXd4jjnA69X26pxVRHTotRD4XPWNoJ2+H9Vae1QYPjmISM8zXz50/rVmpKe
kNHY8bPaANYCVtwzLSJfsjQ1OpZYXfxkGh18if3s96tOvyBCHukSjYjzzV0Q1NrF8vkfkIlycMIu
drEiwYNdGVKTuri1u1UaxAss7R1ns1l4j9pA1aRgBq7pqiH1krQ6cJOQE0IIX2YL+YcWLU/pVnMx
eJoY9zIrQPjaMzokq9Qd6U+4rXJkCt3lcD5nZZ7ydHwCYfI4zOpeECUjndygpjvIGwEf3OKgSoLz
nMq+VqHScB1YH/3GxNZesaV3I+S8/q+ztHpiZWIc7bra/kd/b9cGZlCAFwuORFPM3b8ez40qFBqv
cEPNuzfXMGik3+Wjkczl+6VbwWPn5OApKuOI4ppiHzgfqp8j3/eTlA7cFWcjK9VzWJOuCg/x95nE
24Y0kagZjH2uUo+Hg1ycFqGBP/e2z6ULxY8EATG35VjVeJhJUBtauZc62KwtfMQ2GZ8V7yvAQ5tl
00WkJsmgfdx9Hb4/hm+rO60EkJB6OP0Yd77FxmnmDdVngM1noDPhGDjt6EfkXEt4PeU+2sJvOQ31
ybO419a2t5utfvUh97iryIjBd1Cl6OSY3re8xUfMEug4+kszqVZd5UxlWavK4n8+oo0VmtQJLVhM
InLyUMhMVX1wPRSKlapTr3rOhUvJlZKkw2kh5jVcP7DH+HLN55+ROXlNwyRDaq6PJAwC1ctemjda
FUHVSpS2uNzRUekoxQkcTq+X6eWT6asPTi8qwzHXFlRBF/4kDJ316wEf0BIKCvmadkyLfC8g0QRz
48GrLBcThJ+mnMjKoGldE9KLGGBzrR/BYk/342U5qd9bA5FNZSMKt4udFAk8zQLEzmekoYUHgQvK
2HOekNS0yNnVNKz6QKsjo1DR11fOyC+PVQvIYlfwJSOwENT+JUZIRRKedMDVhK36uUbjzmOuHrMT
fn5gV4PRy58C3FfT6oF5klUvBhBTNfnETO6GTexCrtVxp6SCvkXfteYsPNL5Kjf7nGnOeV0WIT9S
yNk9/AHLfr2/AXdlIgP/gYsJbZWD2lLiZCLDa3LofO58sm4RUik5y098bVMzsXBFmdfinZQJaApz
8yhpz3RB4dlQbBc7S1dG3P5I4ga4bicFnUj1WxONhLNxmplWAoQIp0yTsfS9K5Yk88zKTDgazMyb
07n7M00UTz7VFUeXtWrjqvUaPn8KglMbwgMOE+nSD4+7oyJj9iCSf83mv+sXD4UU90Q9FUnXdJdi
Sk1zIhGdG4IkbcAhrTjTHt7Ypz5q9mUhlyxvwS7kvcxeg9H1neIgMP9b3n+cDdWlNNMbGZuAJc/K
2kPrLht1DKv8Ed5EBtMFmqMTkfrhAkJB/95ak5xDg5HfdKxobMfj5Z2Ffu918+WKLae5vzFfHUVi
+SBi/62q/jt8owNLeaa5kUCWTYTgiNt1xbSB9b5/A/YXvFg7IzROK3yI7bj64NUa4rB+uVgvAW7m
xHfVOLTZkl/ICieyM/zbBNzNVvezQhjleOx0RGMvG/y6G6h/5QYU0q/nSoEE3bDK3ZtXNM5X1g36
UymY0XSKCmtBrmFlEMvUFk8OY5zlTkhYQPyZdi50Pw3prrz2tGksJSEPO6jVSbI9pR7Xsanu/loh
E4zbKEMgocS12aQ1jFwaOma9pz4CaiquAqnQSEhuBKlgWf6M7/BuWyE9tyNcxN93wswhMye15jCH
OJ8JX1/dwFziJVuqJDxRUboJ8CApC6WmypTMrJZBNLK3jIp6VfKLhDMvgHVXbgtgGu+I460046mN
qZVszvyzSFkCFEhUaMjfPeCZOkOda4bxHlJ4U+ZbitHzoPzpY8wIYvwUfY+8+9wRg+uUH3Emm8u8
ObuWPDmtskFUd5Ui1Ap1CwT+6ghcN8BwFGm11RZZOuMs5rqWYB15zxLgsCRTEdAFrU90vtBr5Sve
D0i0w764i89lPPztFdvMtH67EzPa+MnirioK83bP/3VMJnlUNTH+K303s+SONtJi65N/vfGgloLP
Ns7xmVsYzxgvtvPRVOueKjAKkiY0HCmC8DnmW5yXuCSxGzhbAR/wLOCs0YunHeaYSf7dh3Td8qNd
tSWkWCMKMjUrorJbnH1wX7ql9tA/uuGpwKTLQP7wU8zqDafBhLp0o3Qi8OoYDuoS2WBNO00VJYG2
Xo4Wps/96zVm2hgf1NkW7qvjyFQXkT2X5mrSq4y+wm3T1pGcFahL+FMzE+VgDM1e+S7g9ZpmBbwL
5vE6v0NtZ9APPi1RyZauY/G7BcEuhlhOA9x9Uz9twjc+yT3cj5VtJoUXzVGHOoaInGzBGHPeTjKr
mVUFFgu57QNkDvCFW2JIKe63IN/id2li5p0+R2Ko6nY8uRGY2gVql0NqwDExlFDgc3aPYqeaBY5R
tYFZw6cWr2gXIzaY6BO6TfOAyrW1tUuwgqW+XtePTqRDHm1NDb1fkFrZttYktrDUFyVLaaR4OOFQ
357cEYr3Nlb627HCFTwL6nkV2r6BAU5cyuUUA+rKRggZUnpaT8IBlq7eU2onRfpSCWKAxdLdfyoM
zz0yUOyvxw1bXM/wT38BVJtEqBXM7mp23FYpf8m6hp/hq/KXQRzp6k1XbgNKF/bLFJh3Ok4rQOwm
FZftWXT/YySSWD/VLR53fcznJPYs49XuUh0kBTVqDZKieskNAyYK4/UqdVDwS/FDsXk3t7x/+EGZ
Ca/DYSH9ToI3mwSBmVzQ3X0DuPmVSXh9BJASi4DuJUIyHFSLO0eoY7Atcwgff2KVIlgTWDpXSFO1
L0O051XQrXoFF84aWY4+E5/hCzzM1Mv8Daz7tY+EdQ3HQrLZK0zba8oVFNdQcQI/+XOJ3M2DGyKe
J67RA9ynJgaDEppmwFOhoeeZ5xJ6p+/jGXRYREuW0Va7yCZ2zpxPfrcbdWfU1qSX0JMWxFeN2moF
quLMCLivQLvYC51thfppVzGUDC7YC5mLrnsJTa25D3lXqrVV92UXD+F2ddY6uGLb2V1bL2ylPpDh
MEbSYlosFg04yPKi6fiTjCaRktVxzJ3MyEyktiQrhnrKmSHacekCV6Nz4JI0B2fEVJKgRTqYe7Gv
7q5B32KnhdMS30wvXxJlAw4hBY4JkdgxrH5FOogiz+19FI/J3T6snexogYmLEavuMoBAJkQ4cWMt
m4Rg87g2di43llSeMbHlnqO2ugo3DIrkIN6vyXqB88ibnj0/rCAFskPRfHx8HJqZcsp3fH21/3rP
Dua8UgyVPqCVJ2w5KFcDspojv0sNyXeM5Dgfqr0f72g15/eG2EvMtn18NL+/ArEv8gPDeVEiJbN4
1jKVhvBSY1Wa6Zl/UCIGL6ovctgvhIQpahKqCWLDdDVbzxQA3cz/2cmV42nYkH0Ak6TMNZkNawEG
GX6BO8/YMBC1pWpgQMINU7xNoissjnuLmtEgZmr/cG2POuqG/zJ8g0L7aWW0t/8lX9rvbeK/KB5d
R8Nt13JzFJQ/5cn97U/dMh9e68+uho1M6dwDsVXo/aA5Wjg1FQSsBl6ZOCv5TwOyDboioyO4LDFA
FFfAl2oDv3P2SavGzIZdeHcFdidpGtY7vhpkeAcng8MJAk0ZDIHB/9LbViAY2m0hjRycRdJWbDdm
aHh+NKu2XXGaHZD6Dx4iMoG7aAWdssbp03bte0FDlH+BYErtVtnpEVrhGxVSgdZjBrUtynZ1X4H0
in04b0JD+tiKLWXl6CpCJjt8LTlZbB39sQRauTX/XunXvR3899JKNcGB8pa4Z1WqsNoQKy2Zu+rM
zSUMLmFCWpBxXhBhLyyTZATdDJJyST/0Jfx5Vtx/4AhxNxLvJZLaLsebd27La/D71XJpzW1Nmhwy
1vEa/DXn2ZxI011YphiPnVvMAmGtCuSBYrLACYsbagbGMy99FHpTyjWrNtO3dx3DDL6EqU4bcYrP
1wCQoiccAt1AexmV7vnO0Su0p7AwPfuMipvZqmUSn7eLEUb3fqlG/NVpTNThBNHJgdxM+jM3tASR
P/bcEBcZAlkCiCgvXJLspmKwKP9o0rMSZUUjUn5W2uuF6PDklb81dxm5MGckC/9ga1mMmLp0mChS
GLPnITzQxxdI+gOWEe2EWs+a2IZFfliM94ty+HNHXAggmBRJaK1kFeiYJQ3g+6SIFxOJ7HigbbWE
NIH2ccxyJ+Zdp6O/LMB6kwHEKCYT0B7xaDwTcTHlwAaiA7j0ZT6s/IdX9csrnp8JobIYNK8tRNVE
8rY5oQdJX3x+qFdZ9opwZF8H6rMKxDf2p2i1Bj9xDYIMC/rOd1p1CH8SAn1veoTnLwm3ZLoGJ5Xf
lXsAAZsIgRcll55yKmPQriJkkw905XzmjfVSGgNkvjLIha+iXfnfA6FrmpfPkZ7+lP3ouYwiwewE
H6EcbxIn4IwD0DJEHdLhkH14osUZ9kWxW36tUGpHYi+YDHtNFKjmCAvAY7egUzXualTm5acCtmTW
kQycvsnll0FF2IFX96SuNLhJ73cLER58DW0Idusct0OYCQyD6YwN8XSREv/aVKZfpHbFxZlat0kM
QPY+VjwCZx5R1dwkcC7kd10WlVAtd2vPbPF61ds+JTNXz3Dnu1oDPpCRFrOgqmZQsXUkNEvjsYw/
lCCrzCzAoSIGQNZC85rzTqIivJak3bvpwh6U+8rKS2GaaEyqtzaWD1/Yd6hWj8hLNRdJVfj4T7PY
Ky2ltoJ+3gT9q0hl0mSmItttoQYQR240L0neW5JgOLRTeHWm6Y/f7X7JgmSQ8jrYeGrtI5wAHxL7
HIMPTrmdEbZUVJSZQpR3T4PX95UKD1eiA5XmHqWYQKrttbY7ui4ZDuJ/sjOT1DpDtwU9/4UZpJK0
qMZdilQPT3sMIk6c4zsIDem/rHDTKamumHC7WMAfbz1jrpTxDlW9WceFUy4VI7Wgdwi9EpOIqtKU
YX41dLsIMvurESFh0oEfzRJCgUVH1uCgfE52L6Y7qKQG01fXifb3XwL0xNq7I4LtiOP1c5KzCGt5
BEZiKVVz6qSqTj4IST3W9Qv1IMm8iIBTPvb+YZHqXFnQ0dZ5IN8PLdJCMcf8NiHHizXmlsCNe2+s
caFVaIBVxpDZsBC7TRvO3MLDD16gF/D+PAKu5gtR0qbG6T2Gl7wf0X2tNuBvEj0PGCBPGdUH+w8f
hBUQnnu4RDFHMkOpPKRgnQoew2DL7Zy8kaMlI8v7CQvY+bf49Fwi0tEKdv3YsF7G7RjtP7vAIZN4
A5S3kFYceR5IboIlNdCIZHcN4xf75s82MMsyuLupX+WPp/YtGIqq5tDh3ClxNf/0xA3Crpb4yxk5
LgGL/fAeYuar/xG913JnIs/PsSk+cEJ9pVi0NWYPHk6OVhhnWQwQMkcnrK6u9oXETVl8BpLrqRAy
RSyh7RJSBa+0xLDDDtew7nZRQw673rKpn0xurjrkIGgqoHs4IivAjXwoT7ev3B+vzsDfaugocDoi
TmQxh1Ow2gm1jRYFqIyRKUOOcx3KWg/az75h2bRgDATMxNfsDNsohm+kdvfVxtcOpXm/cTzqkoV+
CincLajosK1LNhEnmTJsSvZ5/pMSXwJlLeT2SdDE3A+HQehzs9O3vePZatzfG3n4R5eOb3gFNlCv
FR2ymrb+AT7AdVVnYJTrmxiYdQiFHSbZO+puTFBWxsTCIorW4uYcbF2sLfIRsr7pHam4wtZGm0B4
92ilub5RLvapMLa08BbvCcfxGFilBeL7ERPlfbTpHHgd9YieaRGrVX8hVmJOqpQZ+nODz06NX+b1
jUCG26F5aLhlfh3cgNBIzwip5a976fGch2pmn/YOERPmCrmzXtYoEFwBHFrSdT2gYBgBftd3Z+Pc
xYWx4Gy2kfaYTp8+umIcBYh8mJSQnkgZeINXd7LNq+nf8luiZZYTsOwNmd6t0CGoWzhfTVpbxeAj
OgFlw50pPTYUIi4bSQEmopClFPNwBh7abs9LAL3s2RYFaZ76w05mFdOM7z1JQjOa0RI8/86eMTdu
9xs7Ts3dcaugLFZKF88abm4UY7mjQ5x8pnD7c16fF9bdLgUDCFsRDZV8kRC2oCOUWV0p3V0Qwu94
Dh4CvGe6fpBRFuKOAmE0Zhp4V6QKmx9KPK85aPufyod04j+y7Lqys/57/q+b0/77EfT0Uct3gS5X
4oJxu1Xh9O/38uq1vbfdbCyL6k30GfAzumUASjzkYzjqRn8SwhZfFjhr5bwAM/QHe+bhgqNI6tpu
dwGauwbXB4XGW1pfSRU59potwekt1K0TK5rtF5yzLYiXsTVHrEl3jpjiuUrOID+DVcXseibKteNL
M7QZbibKHkrEiRdKCE9WNlofVLuDFc8UeSuBuxGcN5yIQazOSJ5GGnAtgvd794+KO7iJcLNCOsOL
9nWPhMb+4Pi/ncPtcmn8vzq4+5Ngjb8SnCON+3TyQEIn6K4fCICwjWdQHAsrP8mojIJKqOfmlqNg
FUHrFfG3I6SgXC3NWlWLMnuyoGCHuKZNeoRSRaQfLb65rRozdx67fKjSup82FwixPqXS7SqAxpqJ
dVdeqpMLKcIsNnnWt6hE96W5im7okiiiJJ0J1/AJKtehDdqOyWHDdJ1bAYvdfV+yxTMlDW2kR1MF
yEy15oS2um3sKkHjO3pmaWgkGfCro6LpflqKT0SNFkG+7cF0vGUPsh26+Whvpk+xDdh1swLzW/Yi
3MKERbixtsmdOCOi2P3l96OelH7yrngHu2kFn31hOK/fnArPN0LmJFgWWKhw9gJXMwfCgj0OHK8I
0gP3gHMokbN1ri0plW/qLaTdXo/6E9CWc7aQy4HZw/Orwnn4kWTSgAI2DTfdEwinEcnN9MFMgTmM
4FO43sh2m+WlyncL3GsL3oWTxTwJJpjSz/pKySrULFmWs/ZRCeSz05dRXV5xhhv1Bf83c4tkx4Q0
d28cA6Qj7jNVb4GkCPRFdlebDalAIRbqh6ZXmPnK2ob2ZssBsV79O89DMYFeScMzZy6YUkmmze7j
AjEFdujWohxoVrU/aCWo6tnDrkB1bijF8TqI0NiNkucBOHoSBO/T9dMHX1EGRFBoaqBnJ90TgTte
Jb3Sl9yo2YJO1u3eKJQJ0owStDWe2BmD43CDDD1SnD3vCgM7jFu87Ub0/oXNfSW22aGpBboM0LG7
GNnFv3bg+pohYes814G5lCZFmIAX+zferkoR9TMm7mW95Xxj2YqmBtEr83AKaG7Ipc2EwLXp3oAf
gRTyZlbsWGOO06ly5XfnVV4ydhOvwyykRdEF4+1Uhi0TanTCP9tYN/pLvCCXiZUSk/9fDcEnakxS
nBojWqIFTLmVN6ewIPideKLQOK1YkNYRf6qXVoGq4798k17Y9afnVKwG8LVBImM5r7LAHBLZXFRa
mbcus03kJPI6W4LrfwPimnmY8gZdzcC5vOLP/xlUAwngKvQOeR4EzQYURvH8VJS/h/PwbGi80mIg
trrAHkQHELYebDP2aiz9vqR2xZKqqGtwF8zqf0XKZlZ3nHlEX2ZnwZgMHbMg8hZYzM6tkyo86W1C
FrWJZeUUIKmhv4BKcuRGZo2SCj1E5BXdwjpytqlDotjlqA9lzNV8r1fMJxwwLaW3nAG2HHuL8l8M
2wp5adHlhNei8Ida0D6SmEg4wiaKsxTD9/zS+TngLC5y5YRZnNDboQmxPB6ftr0fgax0UjE7R4cR
2MT/NX6Q2bynYMfUTOfEaHV7HxOb4icJoFehWpC1yUMMYwTWCDOX9wXCrlTNRWDTdpdjoEyLhA6e
9tKHIZGMD1m3AtV/DfPtGmuAPLSdLJ8GGtCb+alQVAkcMmCtET3qLTxnp2w3Rlzon7DLQS4KC+0n
lG9c322nFTVC7H5R2N+DSLdBtkYPtvRG5+2CNeXh7eXBzTJgXZK2bFcvn30v+7RmS1TvKkDD7DPI
tbA4ImuXlFCOGfk+sHHhO54+OI9xeGeDm+1HV3eyVHafr6bqkDVNPYzzbswp36DgFCSOK4X0vHFo
81IK56R28QswvtW8sMx+lf9jfxWZMqLzmuRru06xUrc+X+tq5HuleehOYvQ4DhapwqFW3a4z5LDr
pTSkSQPbsHxCWw0unxR6skCbfDz2cd+uZAaeX8ovjWJSV85v14ZZ0fgrFvgMzRsxPX40L1N4Bhz5
x93XkLDJ4X6YvqpSX9+ugEUm8x5wc062toObqMnIv6rEaxYl1mfyETHLWiG2YseDa1t+I2AoIy3c
ltusKConmHT1mJr3Rc2Vk9MVTB9GRDoBE8KyqmTue62fNqGPNXtHC6q0Xs3wnsxrDRSyntBb/OEf
C4gKga9oAg+au1w6NOHN2Eg9bHmOXL1kk2Jd6aDXGrDTUc1U+y3sMV+1MBCHZ8BvmMo0oP/O0OMg
k31hjI3C0Ru4HDwerSteb7rIYtLCcNqaeQz1yMnnjMrY9AxSTaYEE6CxbdWltkjYM0bQPZRw4dTn
PtQKesALwvueHePH/QJ2TbJ6KJxq78Ey7A+UgCn4CS51D7d+9f5/dN7P6qnc4jobuhX8jp4XwW9K
KIYeZ3eUZxt5CGE7VsqnGJDl6uYFmfW98fDOya40CwzfahbaGHxon/onT5qUFouOqmFF62EyvRRy
szXtF+R1BAO56oUxCqU1CcdtXtyCWNoea7p8zhjPGVjDY5K9fCMCzObrS6nMJ7ly+63m3vWg5NYo
1I51LQmkB5sxlT4kx+hYHzksZVj3v4ZLOnWcN5lYHyPuNWBsXdR3R6riE76NkRhorp+Rv7hRxN+K
3GIuz5SqunyPhjDOd2/Zbf0tEcHb3JB8HU9ZwLebEsAfvHvdOHbG84Bpx85g7xGSwM9PyAScsuXS
QzoXaqSb0AlbKduMHM36ZJPPJS8hOrzBixCRvJlpa/PtjN884Au7z8LgCDalRtQEPpjh88keCJFC
CkYTApQYd0nkb3BxhOi8sVvbscxfWyyKDCd+jTeBRJr7Q7ZD5HnAjX/P4N+p7Vd6aiu/p/8XwePJ
gsZgkdrbqgFcK3B3wRmRyXRP+HVqgjZmslC+GuwBO20RUIuOXs1TNnUV0bGh7bnyfbB5LcZVBNOz
x55Jzab5oMm0cX6TJsZ4/xFOlum3q7kNBnS+FKaoJPjDfL/G/y72M+B7LQXDhb8xs/S8MB9fDdIW
zPVAypwgfGYFdKtiUmN/Ccr6XD0cnNtocGeLL3DvJNIRLzP6isHe5oGza0yR970cH5v54omc2zuV
A8l4BRPVPu82QtMjN/yt77hkdwOuT1iQPqgfYHLmBYELmqRjlk5rPNu5EnPbltmdve/58ncfNgDd
JuV1ewcEVbHF9B6cmROo03JDhnVv7cVH/+QptcYY/PderqPPYMXorsRkOdWzvhHeRg/sdKzW0ghm
eM0IOVfU18zSZo9w4Q4ey3+6qePzsWrwPpQoO0f5ZZmOjl2iL7FdizgjHSplEWZSNaSi5spD3UQw
K0ee2VvVXpm7tvgdpvgaWxIzLCjz53X6KjHOlHx0JBoabzLsXka+edIKmmFkdzoL0bM8mRZy/K95
dc4mXw5k8BWDACVP0TsrJQFxf6kgW1KLHStGR+F5krttljSx/YImcLb1ostIfi1T2aJs8HB29Md6
tzA/dhkmYrGBWpLiZ2U3cpbPZrCOw2z3I6i/BQKv41cjyymOE+h2MJDjGZcg+wZflVghnJI2dKBL
bHlG1ji8dRwoVVbCt/CTNYIedp7lBN8BhFlwLBZA7ZFYTkPVLCNsAZYN7jtBWeCIC5bQ18dvxLby
aICWE//Ud6DKh2n5f13xwN+XjhGQAqTcRh1jYKGROrPHgF8goeBljqM9Mp8aEsFGxlMQmYFygBWJ
QhSSDRd6/KX/5t7gZopbFN33/A7VZjOVNW8a0E4UDH+3HUp4WHzGWHOxUuCw1n1b9/RWBKMyvbsp
HU8bv4YXAEab5ef23FRLvyMYAFTgZdHFkMuNPLDo0LN9oJL3qoU1JyERPfrdo20v4zb/VIALlk6H
1rz28jTQG+WxA8yI63Q7HUQ0J4wp6tl+eIX4mOnvZhx0YcDgVMaPWvCeGsozNuTQLvEi11FRaN4E
Og3RYtkJ6cNp2ZBJ/FLWeoEyVa5HIjQhMw5/mKZpS+k6XAm2NSqBFFY90ACwm3fUvDSsNZi8xiQE
GEDDDkGIwWpS+ILuKyT0QcrqENhUV6CS1vFwQLi+zG2QghZ5I7DKTAbARHhwRAQQMO6JPT4eRqXl
iVMGF8EPA8ZswnhmA5t5kemj+VDrvrvMgiErBxcthtvFs0hLJSaxphEcIw4MftGLrK8Kfwg2iwPV
S9cUuyWLxSnvsHo6HGNM/EVieYiJxAsD/bjoupRvCudbRx4OPgd7D3NjOz+GU1Fvk8uQTsC9xAHe
krVecQk4KBxVh1oS+211zKKcU1iNgmhPZxkV3D/taG2gwFwPnLsSyAKSbeY8wmlDSE4Y59MVOgv5
UtsbVcrhEjxldaXOeVHTuswP3XUKj+iIW/B+R2syDcU/W1ukalGNA1ojRBcr5Qt+aXeWyXHLhllj
fitghzUYeliVZjzlMHzWXyUus3SuQSwbNU5dn39S6bJhFz8zfA3dhe/nz9lzQyA5Qjzx8t8+QV02
75kzJmaJ9a6mU2kITvmEXwqilr+OQ/mO5CXV9Sofc+j292odg0rxp21g1bmjVxs5gQak3WURzijw
4rVS5nVCbTuxfJxcjOCiQVdjt2EWrQ44GjU5/tZ2qPUSdBFkqeVRc5+ZpF4k4lzNhP4UNyGuuj7X
DAShQl07xTzZV6o9M2aJTVp0nfThzRKv/s2Fqe78lTdqBg1mAjlmZ5yy4mUHSXxt6CnZM5m5qhLD
lxhOZO6OEP/eE1BEwNWkMx4oFKXew5kyDoPwBBMSN9PalZcDwhbQS0/vyKO5LIGenkxpAJBQk6+m
yOxidy+ITRdr985egijfaBGcFqixIfBEJSB8lSrst4xbHaSOmG2QouBsWjALwqK+SDm6kb3aYTSk
DKEGhD5iyB/NSAJrs6Hze29NkGjwtR9EpLXVTQJA5nAvhIJnz2QQSxRhvPXSi057pgzBwpD5RAgo
vbka2jrXiEFnPQDRKiq2yHChzCvHG2FUml9BoEcqDmuGHErsU+R0cit5QmsDqteC4ZpuAt1pBfuD
OP3tCjXzpztXWUIR82n/eAu/Vx9P9b7b+rMRA7TyKrXiR7TiQLLGYYgNsgOaJxO51lhfrUqxoddK
zH5oQknmaoS+gU9AQb+vsY58G2pkv6CLjf/vSYcS+ZdjP91ExZxE8ygh6zsvCUD/ravaO1RwRLpy
1UsEK5Y8Pk+vS5nVSmtXBEJgF93KLMll+Bo28/3jjEKXv9uYauGSQksSsHMvMaIavH6So3su+NRz
6lDlLt+7MzMFfevJmP0TIiFZHi0BsoAYRHHIwAV4Tov3hNXavZjJ6ZtfPenqO43G658wmPcYJCYo
vgoPG1eCf26loCnQKHSKXhQuOQ6NjpIRHSf4WeTio1SF0iJuSvFm/HUvUmMMs8mRL9/nz0bMiAHT
/pTe1NVa52w7Fvumb36mjbu0pZxWvUZQJDckx2LcRsnCZALGYwhVq7Z0Spc0/+5TnP2beZp8n/P+
BihbieKxEc6IPkWHW8YAcxNxI0iDL3eLbX3CZR4pi6ZoqqSptBmoOTnNKVryslz7jda5DiophmZg
jcFa7zaomdNeEdusQDFiNs+IjXag+TbsSK1DnZm6YquHWDmwQCiwouiWjJ3DXrbQwlNOXu/U4/br
MsUy+KOb9g9ZDKQWgfAC/0rQM4ZYQtGxq3EAiASBhKoSm+w7a7jL6R5d56qNr3hMObsb0SWcDNKZ
+d6WGt+fSqSAXcjPqgmvNSlAW8b8o3O5aRIJfFLql6xvkQd5SVa7Si+L4b5NRBRC1G0ADbmKKxVL
QnSGsppK/eRgIlaa4DbOv03Dtzs3r5LBPr8yaa7MC+Jk45tgEj3VMl5PS3oDk4XwCRz20S10oAo+
V3vJ7AEVtIt6k1e6jAZQAkI3OgBQVbxoAVUIjm6mrjokdBgC1PKXp17VoN+HvQ3H6KXeEotjz//o
yJj/3V1e5aJLQT95+vH+9T+qtwi12sdto1uSs/qv+V6TJOVSom00cxcLTG9JaUCq4JBugmMp8XpW
FjJcZz+ejE/zPJY/OjF1i0kxOJF+SHcFdbjgGF5ZO721wY/xb3d67C5oYUA3hzJ1yZDjUnMIyi16
qFRE/qkJqWGzlgue3ulwlZqXwDqjqdDr+OnZHxCkZH0p6essZLU7uROTWqTluCjRzkmeITSF2E/T
hJaKG1c1c2qSuVQHkkNmaM/vlTgTfglVustjqKohso2ceeNlOmWa/OwhZmOUtsyEaq1aVvcY2F6t
Ho3Mclcs9+sLQPved0dwMbNI+Z6NP2ebHQ66/EyBB2g0kIVMSEKtx1F2BF7IhJDiz+VC8LxWW/TW
93R+baos7FQ+LUKLffsy3cU0+NrAIvYrStLeifUDZqrT5GL8vyYLi5yob7zuH2Jl+JTRy5sBcexa
FyXqSlev81idIuKH0Fw6upX+2ijEMv/I3XqAfZQ78yQGK782LSjQ86nBmWs6tMvIzsoL6KkP6znn
Wo1YgzucGihRepZVahKYeV1TFBkqMoNOf5kDUn0GjmUJ4ZdaE2jxtV1VtPKIdbdwZJfHaqVY0OX5
0YmoclbEu7GCNfOd8CxKHEj/BXtJA7V1HmfsfYACbircb1tWLZKZeyvTN+WReO/zva6b2DzJiofX
7hiduBy9cHAMRRPPEoRU51fgkzTC5YoDEWQP+diFoDWkn7oIw8osNneDr9j0py14sZ2qtgWjsK7P
39vY1F49lThVxKwRfw1JQx48Lhb3MBeKO/UZ7ALPyZMQTaghhZbOr2zVlQrivVqnYZkK7Sb+FwR8
yKHtMZaAQb9EX9fO7HL33HhPoTjfCNLPpSt5WH0Noe5w/hg1IRT0Le1GYVWCqwH+SU5ab9onyH28
0qDNjM9E8nzPUtaUJmHW7ijj8FXOdtH9cL/aRn7/6MHxZ2ZhFb9uaMiB/Bn7mLLmfXTcYgZQsp3t
H7pxEePEnhvDCyz/vqcxvBA5WpbhJOUjhA0vVuRmRkewyQsgl0Hg+PWoRIvzqTTzf3qundewauHv
iVuDz2sPrGGJfw5autbgEzFfsLh81ArhO1i5jBtBXLTieE8a2V2+DPqYRhoIKVZ6cnvWAW447u0y
MzSGDM7OWwjO2dR2Khkb7XXNTytq52NqM2Bpr0PV3skHRTxBBHO4Ke97p4WgA6z1ZFXS/4hVICii
r2E2VjKfArT6BJ+1t9Y1cxf6RlFhqtBS5C+A67TayAcqRGQQ4xeg4UDUqd89p5aJgUU2srHMdAOs
yUReUECMwGCWdeY19n6sIRhf7W60HPG8Va4rhUaQYvO5m66SVnjt2QF0A+ywOtc03HejeEiMo7IT
noU3/05B+6iGLuxOLxIkggEe8VF2GniKmsTqy3S0Q3u66/F+yT8UnizsmCF6WOstC0TmbShIIIcG
gnG0jaJvnzqUItT2dUr8Z4HykeJ/getUI9DKIHw7jyD4u7DqUQVkrOBPKlrJdEmLYkrL8jSVL2J/
tqf+1u9kkMlhVqoGf6UmZKV92DmOByiD6SW2XmDxx3/LLIHxkwtCgbp95U2ogBKV/3nuudtr6hGW
ICkevNoL1j66fOsQW31cHzS403yBLi0PxxXO7F+uds7DF92Tqfdc6gGHNFgiiFgZsncqJltwt+nw
0ZDV05QW4Nbx7GDPCEqp5CnO+ITCufEyEWp01MeXmQr2qvf4z4iaxzOfQ/q4x/D8NB79x4VN9OpS
mztYsvjAscUT8U96JoGb9qZ55fAMpMb/108ip4InMUoPPHeS1o9ZxEZnCWsyr22wBNiyM49kp4vr
kSeiP5QGr8gTPvoA6QE8Eh71c80AOnyRPzmOy8aSApveTnAXoL8K2JUrZPdUvpUrsALDqfOXAkSZ
ZHCGANpL9+c8/AvWW2DMkRMHGE6T6pmgnOPi6doklKPvSfMGbol5uf4+HSQKLeXv/hQCi8BSl2tr
GVNv3mceuus8ibFo/8f4BT9DK6MVVhO0yGlgsiF6YQAs7xlBzdiG4KJEwxX/QwPZOkk+1HZ21OC7
Q9J89V2Pw+6ytO4bVcG4qy9ZbgDuXfY6cDwD37crkv4fpltJLbfqVUcVVOUqNsGudlkRddpgEBBx
QdvG0U9qxuWTZ3gSHDOvtCc/n2tyEWBAdY2xUVDDJRJPF3h52QTl6AjoLk4Uqf/et2tuPFEhRQ51
ooBZjiFSGKpMNc+BLcThtxyKp7s74jtkvs7z6DXcDO6JTaZadn8TMwEctFsoKXHfApqk2vOGxDNb
tqqHK1UKXWOmkjdVA+bn4nTVIMak4t5U4r1NtIL8ITwFhEVIVB+lxwEpkNdLnVcD4/rbuGQGzPh0
J6BsqZz6aIdKlMH9TWvBrT2J1wQc6tWflSuY2cPnxH/k2MI/QuMRb4GfO+1MHwJFndDLbLY8nlBt
FXMnVjWahfikqRNL8WdQix/gQgx/eIVV7haGplTRgxF05fCcnAo5TILN9QmDPvyHtG/mhIRr7Vif
VjidSAO2GuVpUEOu8VB5GujyNXtmyELg4uIxAlFY9o4V9yL+zRC/12pBmh82kmm553WCCBJbhT61
kY4Xjao/aJXbfOMgr0GQEietYolz369u3d+2U9ERHwXzooZtjVO7s2wRWAgoDflSlZ5gX71PsWQz
oA1J12D4mRJj1J8KSmf7bJ5QkmKRDHvBlvWjriwPJhpJt/99MYJUApmPYxhLl31I28iI2HaqxPvV
yKiEWyrtAOGj6aMIOmv7hZtoH5JqOWo3t69445Ci/q+7sGM/hkDVuYKonM8JESyyORAnMuq08ldn
CbSBPeUPg3n86pDmWyIEAKdeMuWKWHZdXVy9dMXIEBlzoX/tF2M5SWzHbuzEfE7fsRfa9XM073Tn
UUkw+D7c6yaG8Vd5A+wwX7f7u4h38hzyemwwQ758X/d7HzscJhc0QTlW80FzrLXXPho/E/FNE9sR
gTK95rkTe6Z/S4N+4sYGbQBVyHD1ZdpB+kH9XC+ZjUZEPV6DAnBQY5lGfls2qUvY5xvslkm/hu1V
ZdbPOg2OIb56gArRrR6viIc8mrmhPgpECSPyGLHGO812HEZIMwndXsLxk/WZdxXqM5/rDa1tNnPS
qyjMe9lB+ZzkHVFvpifSYS66KVF4MbD6fL0rId2O4oHIaXQfIkq9TmP23WpOfQVceDspXu0ujmt8
C70btkWUFxNkzdFLznjBixFkhX+K7F1PYn6GM79/riAVUH1lQTOnh5gaGQn9vuCtMVQIJ3K1KZl+
uvQQ9iuNswTMfdwWZIv45E+1Q+NCnYlxuT6D9x5Nf/uUy4ZutEq+sijbe8XZmD2cnn7o1o03HRBW
o8vmSW0BldYuD7Pda5oYhtId+/FdkuWsopuZgq9UIKkX9xwMf3MyCsaVZnzz217kTnFWI0Kd8h6M
WQexZMTN2omd9K1mw5QCo4EC7HpYUVCxUzEhIF3fOh2Jmd7b4ITDLhQLoKTlvWJARrKenDEj+ZfS
WDXCnXB3tKgo/gAP1KSx7fQPGoU2vb2h70a5k+ukyhs+ADNZRtkkKRtVEjveteN26+C3kCElDT4n
w6wvxRrTZlhof+haRVGdI/urkhl0NLN2wO/g/4lVDRR9YlaPkeI44YrejFh3garSgl53GcFCcjHj
92sr7nrX9qL1V6OJz966MDoOjqLXZIJ4efIpmIOt9XniPZc9eJFDvJGEwEg7gc1mo+GEE1RrYIAa
ZTu95rHSsH6ClJFfpQ6wxzvkksaaaFVXBLAnYqkUffBZIqosRoqdUNeq9d7z+SNaXowZ5bW8bHpO
yHsCPNLK3r4oolTizVzbXyWvI7FqAQYpkZW1ZSomy2uaacPijQ63ijd6hCwXBgRI9eRwg/FNAP4r
Ni7X8/z0di7+nO35gKFQ/GO+KBze5Be/IzBa2iLAEvmNGez9QIXL5gs7F5jkQ1dXN9I3Brpzv6CM
IZCVZ7TylSWgGaiuyaLQF/K53Tdep5A2LgpYZLUGymLJ2ZZq+JcHTyM4dtQDGulSxRS1rXqmSJ2x
Jh5YODaNORh8ChuHFwLh5Rg0TTjHvTIhqK5AY7qtJhGBSzh5+yuyBiatXSKU6pDAVxvL75GV4Vnu
4TLK5bPK1AzI8U316OQVUngNLW5d2oqbBWKO55cxyTwtis8fnxhP6ueuanJZKKF6ffH/lnnFPPG6
K7doF9JK5TdTscG1M202fYP0QlmILENRL+yzor2PfAOr1rXE+zvU6gtnDpc+N68e0DQ2r7f6wpAE
hDTu8k/dHxiBoOkYOchSqr+NHNVeLRV7hXlYUoEsYXC7MsxJ9D/8NpHU53zwXzZnv8SB/2X3PQor
wzrBoXQLtO5g38deYW+6f6sx3gOCXCZo0u1AS1UGDQazL2i5dS5R4rU8MdyNfvQMUhUkXYen6JN0
SlV833npIyYn/DFYxSSrZunMvcZhy9nm2d9PPxVn37z162K7KRV0R4ciOq2uor4FqsLkKD5p1Sar
wAHtGzGibiqvwMcwxwrf3y1qmMx/r/OIttAXZlNLk6LIfrYQMAxepttNwjowgmmuJMGUlyGTfojq
F/5+IZ7iOgpjO5TVlWr9JykQLEiIEcdVRidtEo0qWukuhc9iFuMpFgNd1d8hmNEweMB7pVsjmvPq
/e//BT1sVXdK4Uw9m0SnxMXKyR1ASiKu4srY0ghZhO7rxWxz89QWCxW3uDZjqIRuEk+PJPY6wKdu
2OboQQ7XFPqlxZpbibcRbmQdMGBeZ8dDFQsYmlvp+uu4dFigHcSJBoOCveTdghjX6KJxt8N6McHE
DaSxEa/G4eRT+/vc4FxJV9pLfjAw1oej7Vh8AGLX10UyKaEBcHtW0pFPOCOz3QyHRGycYsaumLMs
DcBhAz80ZmgjCANhIsqY2dEvP3m6KFp6nwAfYJUeTZI9RVmwrrpnH1zABrl8b4eEX7vyAj9HsQgb
WHx/r/Ve02mUapa029ANxkFiUTbHVPuemdN6SOMScQcd7nlFApeGUhUk88rSsSW2nCt8wDAJr5Tw
/9MtdqnawrevAH07HGSkyoSmOsvgMa9sPEjZ32ZxKz48r99f31X8KAuh0G9m6nrQmPvO0/Uk6R+K
mY3pAjFj9L6L2YyCf6+fbKDOMCmFHx/8gw6Txo0V/+XMJEXxjL/AtUPUvw8kxWCriJnPqUFwpYXq
Sj4Tfvh8yA0w06zRrl7IM7pnuZLBF1n4lg+YJ8TPwojscLoQfA3yXVqSKch2sRrNeT/SHJdHSsW+
h1CFL4ZIdI0ShXOgTGHLfUicvLxJib/4jq8yYi09m+zlcO81hT1eDbkyECxkBQJKOIxE7pnvNzdI
YWRRqWHnYt6v+AVMXUwwLEUxlc6N/cw3siv0jznhRnCZb6d7U328COMoNo3b+uGEHx1tn31xtvlN
5VLa97wU7HW3ZZsrSJnSphpq6Q52Ogq62qQPyBPm/LidOWl9Y6TiFcOiG5O2aDbFOJE6VLT+9ijr
xyy/LrZoFIoDKl/VBfIjV61yTkQtPWZz3Q+HBzf5haFi3/2H1eB482fwFgMdspBoXPi5D7fduvfa
vL/vaBJrifMIpos1yT2zD69QllVtVHyCKHBnrR3oES8BtcuefJ6j7+1WvNkwINKlVJKK84LVptwb
o5S1MDUA5RG9qnWLhR5ChrOYhFnX2zFN/O+1Q+O+kpDKz7rWdxdsJMziFLUuWiCy8opB+5F/TKFU
uTpCDmqJSxsDy2TaYwYlkC4aUmZLfzunDLl0vNuKpL+n40iWEbvqvjNZ3nUVUwBpzkxAbsACGPyO
FaBo0lsYNoUgB8nl2ZfrpdFNB2YOQec5nD7fc60xCt8oiDKX/at3aiuKkW1VtoS6RSiTHRHT++hN
VjtesggHgyeZw6PX1movxiytaxnNBl1cUb0/hPSJFgBA2s9gqTCVwobeeYlgCl+ADoAVvDyzqekE
tJO7wKmYbllmuqLuZgVmC8FcXDMNDF5+BD1klBHAoG5aaUxbSfHLUBFA+Ajx2TWuA2G5pf+Q/Rf7
lUmma8YBiQz+8+1oERt5xhvgG+5tE42d8l86KTZ0Rv99txgMAtJvv5M88r65jRZid57F6hUuAcz7
0PkxmrxLcPO09bAGbrMyO6vgM96PUqmNO+xuHg+PGdK0G5DZuZA1gHt5ox8err6h1LzHJk28RQzC
JLGA5X4QxvckpZBnphodC3NDiqUV10vJdlDIavY3WmWvdXuhCgMM1nHjReMmbjx4DpYJVCJRT8pw
vL5Q7T6lROVVgjPrO+6Le3qo3QBWTOLpFt2wEL69/+PYnLHkki2ljvQjMjGPWtPcojyaLLSeIziA
UeTLEoQB5rlV9vSEPYgQCe9/uc0cB/kpn7ofiQB/7W9kl3hY+Q9MXdM1/H5sFvmaTjotYquO+DDV
zv37yII7iA4F82fEqZumaagM3AOkNfqE1E+djysM6NR0VHfLJQ0LWno4YRZhf4mOiboThIYxOcCh
ZIxup4xG2tAzxNrw8PIyABHw4IaM1SebI3SlYCJRAPuq+v88BQR1dQoC8iDkrxy7WXkuWmWMW6eA
7G6W8KwrMrIv01xJxNxvdjQg897VDTPoGd8NJwkROJXxAnXCcmePyVH5JWrxTIcb4fL3wT9W11ha
fKLoy/QOZr/Cla+KIPhwpoGUcvzIT90+DnUTDUmn5EDKruh13A9VXISsnA8/fBF34O5705ohRPot
VoOrxj5A4gwsxb8H1Tu1898qvXMkCX7AqFx8sJg1rlFNq92miAwbCCnphk8IvFejhD/CCetJE3Q5
bbEZyUDHr3jJAvKffxO6vuxSZZl2ud3oYcgv5GrhC87lW99B26aSvMUrNq5hucBFBwPlNypT/skP
yqh9VnsXR/qr4LN6TYS9x6Qt+Ic1Ik6mqMzVfLpAW4VCMOygsdRwM5/j1vEaKjpAT4q6eQcFKp5A
ESm/apnM05AJbI6+dlahqhyYUbYODBDSyshr/CNzEipcozsIO2ZT96mc216O57Vecm3shqjbX/Dc
QpljijF/D91xYgedNUTkdzPeGrbNuXnyI6j63PSE6+aUXBjXTo65xnKJUTTDXu8MhP4o520AmlYv
NnxlrYsZ8GtiJ/kOhsS31u3nFOMb4lGcBVsN5BAEHPWUlDqPMORFCN8Njlm8eS3BFTp07N1Rgii4
RtBU3bqDxVQftxShvQNE4xMsJKIjNXYWOYSrJsiMJHqH2PD4KfchrMIyodWf/y8DOv52JjA3ccY7
7lVNMIGazUWYYHZDew4ovQBprQwRIVDBV8X3XhAzVjTy/ZIYJWqMt30N/IOSUdgsP7yUOiK1d8Pe
PI80VY7VH3bLcpOOPRMriUYHI9PKzLm2l0eI2mr/V7QkOOXZsT8HAYIa9YqCVROUj8qqkmPFaeN6
Ll76+HkZu7c1eJfyIPjKbATbiKapYKzfcTkrr7wp1TiOI2YObcJRXoEwDiVUigcb/0BLE110+c2O
6CuR5ZS7POlJZvSiVwLxtUqfAaJ5FCi8YspO/lcs2KYFdENjOeYOFqHfiGQXsLC/0CmzH17ZJUrL
LbvKapd9ieLE+MUQFeJ+p5LnXe39b5/dz2pdWnK3Fkj1xklvrQ0cX0fcJtyZWK6aZ5K4LV0w1k2e
90i9o3AMtdwS1yaG+oF73QesIifVF2f/zxW5NncIyqBOLWhLPctu6OZjYaIJvetDxgruVGCj95La
gnSEQDbICcf1exnXJroIJbFOLkx0d1Kfv5aipae4ZejoiPp2mV3XWlKWfD2iM+UbSas40ipRXiti
6tu/QK0SJ9h9xZUdmt8mWHUNSEFPoAj/dB/6wg8R9h2Ki+zs5kYiTojAobQ4JMYwXStgG5hAc6Xe
Q/cVy/OnQOaRVLPTGjeHCj7vUu4vYBPMCOtBMxmgZ86INfq6BcIzmJAOrlCsuiJBEkQjltr5WR12
++1n3OjFuc5y1W0rRr8/ot8di0W9AIDwaIJCdpSvfsnM3NpbmLX1lxcvdaHunnCa2q8Q5z/JoTdy
PqiOwOj3NPfeckBCRbyHlePlIoXoc0w1OkSOcWbcL5YUMKJRUsd5ci9TK1adB47X+9SsTRJ1SHJ4
no7Ftj89Szb8hLCKJpGXtOe4PpMgPFqP7BSF4kDut6GASlv1c9A+L6tYz4JBZcrbZte7fAB5pjOp
Nh3b26ExipZf1HYZPtEJctc2W4OYYDU63PtUMY6N2RH/W4ViHopeyiLI39h4bRr0Ek50Xl89p/99
LMhFNfKJawfIE4j41b9X0u/Zm1r7h4A035vAT+0/1vi31UruVJaynYNIkTN980v8gE9eJwB4O6ky
70QYWFffs0EYG8rmYkiI/IucM5PdwjqTPs1H0LzxsnRtGebexEsHRwhzipSkK6CtmwFWQCvaheIj
3jqIvYCaObaeHxsOIGRdfFyva2dIG4lRLRSlWattiR6/uHnqaTWIGvt5Xd5ze2+rMxdzxpi8otg+
xHw5hXIjR5Zeql7a+dRBD9dKj/JACaGpVRaLSIjJwzviWTANquQbvU4z+bFh8jP3lj4/2KhtcTUZ
hZWLIbI4vYOK76SL4nLWI9fGgSGZytwO0wmoVK2PcP6b08GOro5V2jFYniZbtH0mKoCnr6L+5fMT
Ku3f5LYmRGp4qEhHlOpoGbBauxANN32CayG3HEPSNKnT2hBdlhZ77XfiqYnOdaB8b5fnvXgt8D1D
fzA6Fv6nG55JlxHvs3n94f8wTnhAuQgEvaSD+aSVxBHLgWaP4G92O0RupOO8QIjdFSWBqG/0DQwE
IC65Kjt7YZtxm1PNrVBUl3hCsxpKWVnf7Rvnd8gOu3kVx5v6tXpdSGg3/39mscxNZRHLk39+6aRm
PE/pl4ES7xoS45/G7gw9b4I+4llAC1eIXGAaOb5xEByA+pAfoQI9gazU6K2b5c3x/usu4yAtNj7Y
LUwRTb94baxYScdj3Rc5ZLA03yE3zFDjwUM0Y2gRKa+bXDzgz4iyy2ic0FCb+zCo6yh04biSC9y6
hQAJIFv+Y2QRp5bvPNZj7skN8/PtuIhNv6ZdIpa2oq6URZr3Kc/1P5I1YVZdJgACaHQZRPsxiBut
F5lySpuDF+XwrYt44BGWKI9JJso5mN9gOuXFp+R2B8hT7lb9KRO46SMNGo9j25VVN9p2rj8HIe5K
Gw7CP23GJcG+MgWejX7H70e/D249LWn/u2+fBNtQDvymgqeXwyXlbU4Tn7+lQTIenvwvBDz9BS3S
R2mPBssZ6p30QLu8SARGs7aA3wjGdqaVzXZJggas4k4dZ+Q3U3FQBDQmtlwa+b3Y6fU4cW7FYymq
lQksBayRXB90cU4kvhL37lr1jjxaQC3dzFM/89OKC81Fam3uan8sYiDzjeDdXBQFWC8gm7DFHkaN
mZgRh2KDvxjiX9ww2rqp3KJ+pEPM44MWhN/6P5TT+qO9FxF9GIOXNkPzJz3FMlYaOjRg6Vwpc4i9
8L843RHDJK5ml6b5OrhtNxBh3Fp2K4akDxujQNF1TjKULiyK3V5gpgtNHpAo9JAjsco/BGf9b5bx
qV2AnEYyLkkaraG7+deO7SMguvO5NgFom8x5U90EmZV23tEvj2aZCde9G4Bm/YWPndDlamQOIQIU
3Dkrz3A83R/9O3Jg3Q8rS8hSW4mfOSy3iWLxpgZCiXhQxOVdaxoUqEpctYzEjcpqhrEADEnyAZL8
fVUtub6JZpLL7KMQ6Tn9acWgbZYOr8vb1IIuIXBIXzKnMKXaPcrZaBf3ovwh/dMvPbfbi1VRyxpb
UtmDF/fvOoNaJZU3K56g8h90Mi5TyEoIEE9dSCsYt7qCQbcjdhBAmi80OjRhVrC1OrKfM3SJAoIb
Z/8nHsaFK8HCEj+22y5ZEa9XFcKRRy7abviCqOnQagbKKyHokLkD/PPgHgwKdmPq4Q9UZhyLY9ej
WagC4hMtQ81DIltcnSQPfI0OvTojB682+yO+wuPGEyQzdv28kP6KEc2ZopgnvdRxYl1ZkOlx/259
6GqNnpaONgexy8bK+8Tba7aiYQDjzNyqSyWj3hEenbg0HSRzd/mu0eK3Ngbp1UnwWgZPiyrkTfo4
N0JxlnpRu2USMd9t/uDQ5vnePjECqysTugJBKxszmGwBaDU/sskvbuZfqTQgaK/70+pSDsbco46h
56WpiREsmESNrR7Gw9KC3G+NLpAFOnukpvZ2NXZEcexZiS3Cm+wo2qb+WfUL/fELbY+D2x2u4+4k
P87A+PeVfErM5fYGJNxk4/cOE5T3v1biSycXi/T6cdFi2lSB2kJzooaRnk0YnPGx8Z/yGEYBwgtb
nx22TZkvW9eReCFHvzBX/zGMqzrW6h7mkKzX2niVeH6EB6EtZA3rPOIxywfnXpr7lKtVcMlwgjul
yScXW87yXxXTnNbJUxGoKxT2QHwwPWxGedfkQMns9UTvgX04YGs1kNcTZ/XH90BEnVLK8BbXpYQR
FeUX2yTxj74QX70ZC1iX5t4OLhLEHod+BvyYUzr48pptUyhIMqLqYlPwo6ICAuFc/LTs+fHrzv4U
JgfOkhCkd6m27DopMkIMwR2L8qohmo5ZP1Lb96P3A6XuRr9VZGDh/jxlQ2V93iT6/BfpDEiQ1U4m
TG4AUOXjuRtAUQGiju79VaNu1OeiyaLiZKBBkSM+5riWUKg4sxUBvnyCgAlhlj2r0nzgvdmZupzD
GUcvOSIXPK/4/4OVXp1EHdjTRP7ljOa6sJ5r0Dip8w9bAeqL1RuzaCHtnPVPK0ZxdtmTGwBM4I0a
lB4QsQbI6kCgH7/Qc6z35untlyGSOF5WiIrKjexekPr+Ltna8p01wzxT//xicAQ0JGh1ySWcI0LU
z6kBcCijdgflQii+DRsQku+F6GWimHn8mp+lxxmmUXrLS4keh6aMbfMHPbBkX0Imw6HFycNrJRfH
aiTxe/BGcOSnCAvozL6HK9Dqs0bfqPgOxCzg19LgAxdz09rbhPEwaW7FJlj+frw0v00nLm4AdXr6
uwugGxyg0bxCUU/ilXVeNQzIy75iFGKoz4+VTd3ZdAL94WRG9a1N0e2MAeugci1p+D8luTElRD4c
ZYg5SYaCJMmEGW9u6FclOmu/sW8w2CEebfTsGtIuCQRPJ/X5rQ8EHt/cIZBiwzkS/9JD3wjm0yn8
+ktkvHuVTuR5v1R67hNE+2Qu1TuFwuDEd8E1htTY3Wm3Gde0nOimg0+zT+2SkQO3UQWzN+YkUPRK
0J6kcd8NoGgl6zRKuyyYVcgtNpbIjJS6T+F9ckroaZZJKD3zXoP26eZs2b+TD1jtCXKpDOP9pVNv
UvJ2pvwljGha1/76AABYydf5eC2btgYv+ceqeDYYelGBtUjLSPbj2QKzo9PvAcyjZvrwsPxYr6rt
naSKEoEXObqCyu+SJwtccJVqyl+LUAVLrjGK83bbAl/wJ3oNG0yM+pbb0K/1jHckm9eb4l3gwZO9
fPjQTsP+/CjzIcnzqA/3bPlH7rxlmPAyZbVN4AakJ6hE8ONet2bUjjvJCfinyFHgKuqwNb5RpZzU
qF57eKwC583VMZVpmpkhiXKYiOmpFzIu94qysAtKSSKvlr0bmFDlSgEaCiL95NAo6sA55siJlAUq
guyisLWdUP01DCZZHCnfy5rs+AY8Ac1clH3ZXpA1m7gwkIW9y3YlZfOukKsWZkLEhGognYrhhpT+
BWO7IzEEUtbMQqo5imuxAZ15g5dR0nvsUv2Nq8Qf9ssROCALSsNbtqZrhWpQAfrcTX212D1DHDw9
TeclNPJBipft2OzJv06DTvbHaBgSbrsWWF1q85fOAelCBeLKxmKYNqw4jxqfn5N3AzStYwg9a7uQ
lB4ErP43SUJVSa2+l8hutR2rUMclAO7ADRIaKi3Ks+Nk3ME/EnIP1xu09IsfN1sw881xHhFJc5IM
UGmQRZS2u6Lwuvp8W90OiohXPEeiPQIGV2vILMky6UrI2PZfCRkyqH4JjKiI75i3dwC06cbNk/aE
JehnAJDwPcwp6WxDxYWea4zBYGvWOSRBvm9uqVEWzczRAmbAhL2vvh01GeIIIWS7m987wjapqpva
BkycvpyG3jR3judrTig3GZuGHPRgb87Ep9hYFNeTvPwIMnl2auNyzb/lXHrbO1BENVzpMynYX6Dm
JgFqBMsIaLy+QIAwnEVvjqEI7CsXOHcu5mKJ2VohLC2tq/KVXyZ+K18vtSixI9nEHR4diF2tq2rd
KOT7JJ+jd3jduAxHqEMVHS6V9k62LWs0xKlPmJwIuTH/WbQNYrj5wVmv0PUGG24e37f43M6ByAda
84q1X8fhN8tWYffq29csT3nsKArjN7RVVtEVqPIL5FtPs4h2UY8zF71o2pGjohCxdRP22zbROw99
TC5SuP4KP6g9F0ev7Bn5dj06OvqNTr46PipFw3RVT9NBVFJtHGRmAfvzFeuoQmwh5nDeffazeM3/
ZnrAtOAJ9MGRYe4tEBjgu1q1rzyX03KsMhgTvE8ppgO75zdPdmO8E8LWriMW66ntJqwU4IBswPio
Nipp1HasFMGlzTeYXVOosrATXWRk6/0WH2bqldBQ9ii94hiZQZRLG/BEaI4m3vvQNDN/Z+odLXe/
Sn5v24ZlLwcXJ9UHB1CqMec2mlJuKPB70QZrY1vtmXfhwOr1Zk8VNqZowzSwA1H5sTfcvHmxXKve
UnFTZcaoWMlJ1yJb4z5DcH+vHofZIIctB4b7gFJoosKrtVOAYtzyWOi19QIA+MzLUAookOl4WR5u
SfjKfTnKRq0aaA4g7ssCemgfIq8/81gdrTOO+6eQYx2AuCQ6Juyr9EhJl3sdiyLhNh4Rpi2AcK6P
/ut+xUp9EMiOs5nV1A31GaGFXH4e/vXhztvGC5YPBsAgnc571Qb/foxX3+uXb+XdZ8PnytwgogBZ
Hc3s6DmCQt9eDg7rEdxXqQH0vWLGXGGzIY+6dmSpgUt9SE4ia2Sn/XM9ZE3J8ikDnV4u7HECwoV9
dHNSpE2ydZSyxpOY+Age6HjjQTTQnSKjuwp2NZW1yqNNYah6V4HpjGtIM06XhrKr9JlJx0uzFxY3
ofIBJz1BjrBhAo5dW2LmXNgc8hUST8L/jKyHIR4mVBvZBtiVw8JAENiUlRnFkl6wCs4p0mLRcMvU
sZgdquwW9vpFZJyzndAQKdO0PNi1mNSs+huY4CAMm+/gMe/kPAsxFKy9HCJsmM+qik5wC6c3dAAI
9AQIuEvWB94ylWBbtWuFs46SCm6CDahyYPrw7zLkdgm9sHl5UwAKobCcSPC0q6Xs4BhXpcOYL5t1
Djtd0kBqIRP6fRv2e5+UamED9HGVCkDjIwk4376gOajPSLAcgfBWlrv3j/fQ1yNSoBL4lVK3q0K4
UOd/Qq+FsppjJGgUWkolhGXZXBfOObuJw00qQSTrrIx4VTUwbsPewwPc0XD5duD2ZpMBV7AvfMap
6Q3XvCiX5u4kRoO4ZZcsDq3RWkJgJykh7lcmfBCXipSBgHRuKCgi0uOUuskO6w7eHnQ9RfUjOt68
DCuEHG5A4vTF9tHZoYGwnniYUvjbPq9JYtwzbQa5WOZ1zSv+S540jWxJKDEt7dWP1s1bAPd1MQzd
XfI0xTkSLDgtqStip932xtmpf1ilkE4vo5jn4f3C/KNSVWe8Oq8+Vd1zp8Ok6GlkUkFQRIJOCmfo
txzqRj8Jo7EY06EDlXsNBOrHslNdL2W442i8Ffp9IjER/G9Fl7Eh+VQJECwf35k77kGVQxRHOO9S
LvCV1d/K/dRXr4tQrH6w4ZD1hjdLAEB4j+yMxxBLEj09MIE4wlbyt/rbldLxQwdo+rwVlQ6TtIH8
/RqjwYwfQY1p941AwZhFzkf2RRaNyTYS5aA2rFRCNsQRbzoL3JKJUkiqOc4JpnExDPhZVPgHeCNW
3+PThAUeRnNgvCdC65/bSv30O7ymr/vLgd232mvvzYx7pU9LRiXCJXo3mUjRIAY/MMfD6fo369W+
XzabB5RzZ9MFSvArSsEK6bwGPj/uIXkvY7mepKtMNz0QXcIH+rum7rwnVZy+zvPZmwJz16vfmyBf
6NAj1CEqXv98vhFKCSUrKZqadgruSCfBYw4BPOmFcV1uEKgRanuPwn9qGUlViFyfg7zGSs4fy6WF
E3BPscPjljDWyQEt0yHf1E+t6aCahc+Lod2sRnG4G/OplH+fWZXl0sUJY89zPSiXrOt0EXWNh6M5
e+YsB07yDAKLLYyyEfHM1CPXDG0sh/XOFw4qjhnQqbr3wuNYPzag4xIJbwP9cdCrg+XKS00zpAI9
PzdGB7QNTKcfTlDZRplzgnmn+g2GjMct5c5Ju0T69S+MihssCEMosvz5WSzb/5QciMF9/yX188aI
7fyaa57R4GgTJDNOcs6PXDrdRCqFlRuNl1gsfx6A9dpJHwVC4GXav9hBSwBoa7rrWElYV6SzN2Fi
E0QfCrY+dvNwugrG2v+0Jh8kaeumc3FEIxDZMhLV+uFWLyCVO8gGENxqneNYXv3YmyoYKsw4/l66
4ssotKcmX467ylX9QCQJZNSuf+FvG44L24iFOi7o4dLF1sv61LSv+Ju0EI6d1Je9a0abCEO2iQo8
7HxciHagfMeSv+kDC8GbIma6hW7d5TqBskkKhgij/eSX5J1PYjoy2beBrgznbISDx3stqrexfdK8
O7Cy0vBNwmZYZvbwnD4ftRGIE0m3r2hEsRBIf2L1/7COfIdASOxawnueTZymLeivJV1tdiNIxfd0
fbOQ1GzGufcbuMbp4GTnWziBYuvXQiU/U3jlSzVWro2IBw7jbHIDsN/rkN/75jggEcp1+b5s6Pmh
0LjsSQlQal4b3Uho2ewzv/kx6S2U6VIoOJSWbHfDz13ADYls03F6Ff3tGNCBpcoegiBzOC8jgKjB
HKdZeUmyjlrequPkZ0JMqa5CLJf7K1EqOyjBs4cnUaAq+ugZteo7sQdeBvs2diRq9qMzmsoZSf79
IOZSYMkGB+0aq3XCiPyRqXMJqNXkZ0LnrNFXOGtf3OSHoT/QIqqUmj8/wRTe0WmkkGTtKGrOa17l
meI/CI8jdn8rKeBWA78ljbcIp1RFUH8lc6jcQxIVqwl/PPyqidHTBnixtKcevS+f8Ns/1dxuvOVs
1yaEJTXng4aq85xdyo2xaeQC4gIX1pjKLNvuKeI5v9C/zI/bh0w3SbRC3WkAd7Vt9TmbAFWpE+Tp
zik8U7MS1FbnWtu8CFs9nIx1VxdJQ/7JKeLDHSysJ91ekF5J2N234GYIV1yQTWEHlHTkdIE2ZOya
HWq8bhOhSKzwBmo26/ANR8G3O5zNDikcyMpYS/vH00VIPdfOaurDqVSfuQ8+Fs2sXl8B1V5uAXFp
6qhFeQm+kZg84WVrGLLcr976SUZQ3BDiiPQ9fi1/RYyR4ZPsQercz/Xx2xTFeHTDGrs4i5FSkXEA
d+2pMi+Wy2KkN8YzsDwiLsdWt5OHmSS2jo2ipiKUSb290dguQex4hSanmjQwTM3ENjiS+HFEIG5y
x/JbaCorZCYXEahAsGR1wkaaJCh7SktwdG2Br3vfXrTNBKSQonVTm3u0HUH8GMVG1NVyQ1fii/+L
yn5QNRHEidEvix/c40cnX4Ff2WgOMD4NdoircSti4K6vqz/sTsnzw1vzExYTr7sBPmz4DsCN97+f
MmBGH+VnVKnyTGAN7ehk2sv683wtRCdW8a2Roxvddt6qIGLvE6SCCRsEtm7aDKgvBJe4QPP4dcUg
n30WNkVAK8j5ooiK4JADYdvvPGs74awdKm0ed+ZmsjTFQj37pBJ2jdXSuUslCRZKlpY/swDKoqqr
/Nyw4t1d3+yP0qZ3KWdZr/33owIajLlAzahrp1+6ts/bVB5UrEhfWNGSMCgKgzCIt+4L6wJGeGIj
goXp6XX+J2i+JJHsqqB01RUCHdbiJYXER+sX83o4NZW7lQI7HjsfBb/LCk1yiKEo3CDeEqR7Ll5k
YUSUV8HasR6v7XD22fVK90yaET0PXnZ1UQbX7USYB6F9xETmGB2U2g/yDWTfX6UWss3BKynPqoGx
naJVgXC3GyRFo65tRB0SqAIrEk2uSRu5TiGL5UW7dzcaDHX1USnswTxumLfnkwwtaoBNZIN42FLc
ehrXmeO64oRXS/0Ox6Usw2y3nPM4OScahBZZO0Qf7+gocWOnaK8UsULcLl9L+Hm6MRXz+VSrZD5/
zLxBUW6KalOAONDC51njqPJnDvp7i71PMs27HjpHfbX9rqf7CJJvrLcYGsd8ivrEwAFTeV16rbno
du1At+Dr/uZ6gTnPTRPdwK9sR+dGt8jq7u/cRMTmVFtQsgvZECU5+A+43JPmCckMlkjmdOQMl/fW
Tpxo8b6uXzCiGKsQl1yvnqHa0yXSUDfS+CDk/dOGaEIRFI6RVB7AI2vv/HJz/hs1RD3U2FgX8lT4
a0vtSrmD53gLgnevOVishnAkhfiykqMQ5eOu+iUiWWQLNz8x9Smnpm/LdxBrIc6i4nRipiCq/CXP
Vx+Ev74Oiti2SBGjR8vMCerCfX8ODFp4KQGDJGOEjOZT4QkiKmqJ5E397djn5XkhYjNw2cRGrLRW
0eOb1fmtpGZww9Rklf3fHC+RIpnkx67SF5n0spJ71nFndsAF43TXXH+dJ8Z3arvEWqcphaDgecNK
zhiNDnmCwsh/4QVV2YsMI8UDxu1ZO2n9h5RVz42qMokHvBLV7hjUJn4NjgOC3i1FZ3t/ytG9Diyq
2Lhw5YJxBJooSVdSB47AtLIoh/fduoHN4mEQ9kcncCchsd5qwtkh79hmYkRS7sfyKtOuedv25SKJ
BEUYO81Xa2w5sbFE08fWsL7Q3EV1+mdzfyQ3YEcUWiO3wVKL5qocbr4mRxsVNPM6SLM7or7TQsRh
MP4fsXEpBGJ3OSYekDBEVwpJUNlQzJFbOpeUljSZAzpS5qkuwOzPXuIBoXp53GT5HZSpd2/4H+gv
eNgV0GMdi0qK5HvKpbJ8AhuCxXrrjLOmdQlI6LBgD1dj3skHIR6SJFf56adSq2z6PQF5ZdpR7czL
lKAIdLV61wAyqP35Rd94Szy5O+735KBa5OZEM/D80fnnz46cj+f7bV8S+q6yOnwH/cdieAmMpcNt
zHALshoyBYWqXDDcowaD9DuzX3+EKRf8/4EQd6iYJZjIZBxz4THRAMU73iqzi2ag5vS4MGDE5DBy
K8FFtFvxjXroC1DWJnvYSLx55ax8iq1dMeANd3iWdl5ihVr8LZc+zP4NUYT8/rZZao6HI6f/6EJN
RjlSQJcPWEhNOLnljV1yhCzzB1X49/FEpneTqjpwpw/v0U9qjcRe0so1LUtRsShpCmHMqQmQOsO4
1i9cFmbOPgqFKBdUChcYWOxakOQj6IYP5Rdk3dzzi7ae3hZkGoc5DY+Rcp9gC3oyosHrJK8Lt+CK
ytXhaRyfbKclZKmv/Ikm+ly4Iaku/0CjLId3cW4fGTu2yqiKcA4YZbMD7u8vhKLHqs4ncIlBuPBy
BSJRKxYimvEzmo9GGgK1bOAIwzO487MSJuECwIATo5VCd3TJ+RjcYusi8JX14haMKabIVo1WVO8N
dZx6BnyKq/AVSBh7e85LRLrdE3aJUvaj24faoCOxT9AsL5/m6NrXV3xlXfxJHsdm7kZghypFi6Uu
F5U+c5Fp6vHJ3Y64DaSUQUDL9gG4kp/fqtDbJplpbarg7oCKVgVjXRhCSHe5wdyzGEmylI42K73V
X9qUMgJn2oWp3kop2cFaoCEhzgCDKDcR296Uh2Jy2pMFpdrWTdaeNtwsHn/I8ZABqjnqadH+vRwF
KvlKSukhhDoeOevooAmGlTGulwDeuNB+T5E3ijg2XGW8Z35VG1PATQsawH9zF4yYqaZbq5ZTJuqj
ETOszGStrRizVVzf/yPqgIOuztM91XLA8GxQE96BZlBnkwf22IGbfzzDMyYWmAx6R61g7O+Gkk1i
3LGs4aNRCQdrrLEXofo58PI5cXwUvfLTYI0RvwN0ttCypzaDN574B5KqoOmvdPC/cRGeiJUluhwD
kDF3VONQ/AHvM1AGNX15bo6KiBelaLvUnqT/ZweM1nlSWY1uIos9RBUR6V6kSW+6kylz3XdEkv1r
iqr8Tm+IjQGUg5NtQWQKSvSp+kvuvwDz3yUrM10462rEqqdd2qwTrlDEe2df1o/FeK1pF23PivXG
VP7JOgtjZaFzDegAog6DglCgYgN6fLLtMCLRSjxMTz+aZdoUn0sR0SiYJr6punQ5mFbE3rWB6cLW
cR/Dxwn9VCvKVK767EOjpWscO3gYcWKqIIRt5owazOsWaBwvejvEQi0LXN5zPEo+58tnxPzDRld2
mCbAXIfL49C1vnIUtcQ53LqofUUhDsZOOColmkv/kRgZuqR637jIkxMi3ou+o6eICfEHdZX48HLD
YAsWneRpIs64rBMlcyGivHE/cuQfrIj3xVrh4Ez2WGsGDiUm4oFdgakI2Vyi5TjtSnMxUrOwB7RY
bAp+eIRT6ELiVvKsQEfd+CSGmP8/Kx4nbHKr1wGiL4Mqr8gXkrwuUyWs2p+iz/91FAB5VSVHyFB2
CXnMZ3FRPvBtHZwszNYSoV7ITq7uTjc291+DaPI4ZVLOQPmd7YZjNwxB/521PoWGI5FbqaJcN7Vm
D00rVxcLhTnTgqR19ntHPYcC8421bZowhdhkUk8azyTQ3ocZKOxqJDHTNC62GP8gix5yfTEnDkiH
u9BH2maLLL5Z8hBJTb3G7DGXrN1SloT4Q1HqQXfFVEKFrT6F7wEZKwiM7fgqT6QGylbB8YxfZ95/
yoyOi7srPFO+huwd+2PVWyjBMzEnKw8Ebv+ySACKOmgF+XulJEs9cgzHS2++a3mzPoHL1EJprO91
6rqnI0k9rEaD52fa0PHH34E23OByRfZA1HR+fHoHrJAg8Ga87swZ3r6ERYPXPO1ofcMCFnr/dmR6
wZyRREFcDIfHJ8GLOm/Q2piFBleQbGZbkor0165BbSZRlVGN5qJbzvJt7t+DheAxuUP0W1As/S7Z
acCwT0jkCO85ENlSrYXA/SAs82n08TOSgd2ze7Hy2qYcRlFDoKTv/L0jqYWFeijxIETCdXWRO74M
UQ5f7T2nuyHCz1juDYiMjSpXKPM35WJvGm8TDlD6tPdmTFYVnHgZ2m+uLIjfsKX9ffn/A2gdWkDv
l7VMAX9lhYWxhDQBRGl9Cvj7Jzu7cH+yddKSW5l8gcfa/TF8fbzhKmmHoHTKoiEy87VRfJzg677a
LvVT2+AX5/XEunNkaupnQ042YRbfGeIejNcXlT1kxtYzk6zGEmGjJA6wPAeJVg4SSY2Izj/md1pR
aZFd8NWq+pU8f9mlxyQwwwxqWe0UFWd8TzBttpSGDkHHT4HjCkUPh/s9GICYOjOPp6+69CCT7vae
pSy2HRHEcHGRIVsDam/i5htirmHEEybrT16Begsh74tjvr7w053P/yahOPm/6MISvEYMg6/JBxBX
Xn5wEWeejkGJf/FNCcUhfuodcOPftHXzhIBI5c9Wt/tEKoR/+KWZBLUy5SJLGjCD7QZmTLhsH3oj
fIlWu/zBUw1E/jgMRb4Vw7Volkc2+NxYT1Z9OpDJKxgetXqlsrexP+QN5V8WZCF7t4O2dmJk+yt2
LZLWzL5OGbZHMnXNb4eCFx4fFNAm896Ox/7xtxVMqZ4aat6B3dlDcDcQKEMDIi/DM7EaC1tvgSRO
giHnB+zAeyI/IxNnGuHRZdF62FbOMYWo9kYJJ3+J9kKRhltdjNRNvULNH2/DVi5YCQXvwVER9Kuh
tch5m6Cmml3D3lq/sdY+n1kYbSyR8RS0J4yEieqVJL60EWREAe1bBIyE6Wl0lYhJ025RYdh3gr1Q
l3uX3oMpAqN6SiM5FxEHUzufWoP6cmIpnr04auoagsEmUv2tnheQSwsGUA/69OapgTTgaYiAzekg
3Fqr0mftXiJpe2+ObQIkmnsLn2ovOQpvPfxgvRMGh4l84Lphtlm7PjjiCtGqjd2Oo+dsTDF8fnvN
zKSOz0JRIlseT92tsCLFa0oXRbdOPxU54OXPkZWN2ZehblAgqwpL/895ash/VR8QczzPjzJu6Y3t
IV7R3Zm3QkYG1y3YM6ieqirT1G0gg6ESa2srMPFn6F67eqjRyPjOs5BwTHQOsOd7D655hQee8Oqv
zKQh3AYedUMz+7EETqhmqa+DfxZ/YVD1yVpiLAaL7iDfARjSB5ELUX0VQlhmmteA8QaqxSPQyTBM
MUfpDpVbfxx7V6dpwR6fpONVTCz+QaKP6Dq2+7rYDeeHhFQA7q1oObzJtWmpQHkYO1cBoaHnsurj
u4VaioKgt4xxIFOSK3CO7HHNoDSA5TEPlYO/mVufkMpEOztTDm7ojEScnmBa55W6/4szIkKNUOC/
zv6RuR0OFjOEjpA/UzvRTy5w1tbZUQ2JulN+8RiTB335K2TnQBcqcEHUm12gM0fnO5lY0zA6mW7Y
4I+WEE/XFEdo2qhoQWN4FDpYWqwF329+Wm5NSETnnFO2wgjeTW194BBJeib04jUg9Al63EaYk+A7
r0wr7vywLrGQdQdNHKGZhHGEksY/n/T3pECgYXarF4nfr1XyPOhZrCXnaRGT4AlpgKfeSuJuqZlA
K7Cj0ipE1d7FeqGODsPFdyZx6nE5XcV7E2SKUAUv9JUAuuAmM1tG0hXeyHnV6uRz2mamE5QaApGv
htHFA+YrSarp/pNACV7lQt3sDbNPkddQ3whXIJKGhHfLdQpNyONEObceU1Ea/kM4ZblShHBaOsYy
0r1dGmDXpXslRY+RjgFOpSGFa8y20iJU7Dm+Z65oTb98ff9/wjWg1ijJl3u8PVKXcZViXsOT78Kk
45d5rsuoO3mryiWjhA3zpKGG2AcL+Pp1f2/zkS6fzfHcMzJgxAIfWDbru7w/y9yjAi39aGUtemBy
lV7jHl56LY9d067np54J3cvPPu8+pbzBLbyAZbGPTrYArm12l6gYOx/bWRWB+uWHjlXN6VeQj9O4
tzORL/myVko+z2iUPVZDJbtp+8pEd4cm5LBwQR0CL1TKoZ1Kn+8ggOPJ4aJkfzlEr4nXIGjioQX7
Y7YrtspGCIz1502rtVT1+qFRuoGaaZMPOzo4/wCHB9o5R99fIwnzBY2Bd6Yxv8HAy1YI6ZSdyHWs
exFiIE8Ji9ZF4+XvxXuG6Ag1u1muVdwIqM6Dr07LbyamQYUdUL6FYemx3Lw6V8mjD8ZRbMILENlW
GUFgSVAwvek4muJajTzlhKPfyble/9VuBBzZp0HvRcuYEt5mJNb1Iv4DpffsfkyBAclKzzs6/jS3
Oe2lK/Qi53Dcz3XfJoVsXWf5MLqFRfl+fo6wjKgJTtNyT5t7t6hH6Als3MfynALjP4suqkvurr9i
X4tnza16Z3mxiLqEwHdQxehVE/UYVnIRjvChbz0fOdhqhS56cbKVJveu/nujjtPqpnCR6iFqUQNE
UburGGv/BUk+zhR6RqVU234F70lPFi0jhIupDTZJ+16ZQV0amza/lVKl/+/4iP18URL824Gq0hjh
X7jXDrLYClqyEW8BnSJE7DrN7411hz+1EGZN8k9pWW0dMSRy1aJ3UUSrZk45FXUtyS3xnoO6ZLfe
41eHdl5wYoES+0en05WRfOoSpiv/6N2lN6YtFsia10m78h3DcgAIt4q3w/J9M93xqAOPngk6brtV
ckIz1jSgr5K+0YIJb+++LC3SRK9++/3VyN4zZBroUYIAHxN8yvs7xRHdbYhVBGjRH4n9Mr6+aROd
Y8EkmbQ3psS42VC7WCtyRa1AtwPuHExGo6XoILJJVGzNYXrpwi68iGu1KJftv4Ab9zQgddP8ROI2
PMgmyDruPx+32oAHWO4eEOOFeVcA5/bqGOtIdrBhZN0+yJ8BxKtF52mGlxBzN8+9/vBSuw4/JRfo
Tth7snIYWQv4xDVKF/PIGHVv7vU0xGjA7a+JkEMswYKZ9OcMnHJMkBv5OHRZ3v+Mb0r2ZqI0IUsS
5AmZ2eU/gCL7re7vAmqBwCZv7BHw/f/GQi7pf3Y45qrIykolXDGpBt0aMTnQ0jDrGgZAKEK4JOnV
9fsHwDSXiTJkeZD3eCXGrSbx4ctO1Z/fuJWZQPW9K7Mz/OKWFICWut+tMEjRIhxQQ9FzSYQGdC0B
3FlfwFTu2Xh5aAISHkteTuWucw4w6E7VfdCJNkQXmFbfWvD+aABYxEBJKH5BRx8m8x4PfqaXbKF/
lMgHqyMMiAviIFlLKzanSFw23xkpq+XJRvC6KRkH6OCisgwxfLC/IdnPFHwOVFrZboqcdQoWo31c
RvnUs0/CAUCLUX/et51rSfRkr/661LsMmGU9TTEtAxhNY4f82DiWaFqqv6ymOBuJ/VZjTBtg4gr/
cMNc6R92uSQ6pprOZLcMWElTVlNBs5wyrPCD0CeYUkJjpmnuiWARY5y/rl5Cbb42m6GKzw6JQF5S
OikQHwTvzvrLQAK1E+DoBOnHpiz/MFyV1ysbJeX0RPSJ110sfeYptqQ80/zsVHsOuwfzpMQSkIHn
G+xHZ9EKObvPxI0M08MQpBqv2Pog7FHxT3egH/dlQClMxyJJa0JhO8CrUPP4O271mO6p+rhnp30g
7SX3bQk1YXbg4N+FABw2mv/Z4h0ynBQd52WS9VqP0aEs/y2lidrqVe+dRn4xUQ5oQ6OV4D/ngwww
smYufzO/t2UVtc4vOy0KGe0SguhZI9hl03N/1oDZ1wlcwhU2wtinA/NddSIc8QJEXY8JjQ2G9b/E
AzCWaSM14VY4PkYyGfRssjhOjJrsKXuHbTPpCZfT3WHnaANOxKNGpRIh96548TobRcHqqJvzig40
ddQ89WuN6UmPaSgAgg3WtdZ9BDAV1xiO+uOamDUjWiMvKImTGKyk/TXspfJJ2+QcFQHqO5rbhm8k
SdabX4CsC/zLfbMyCT7YN0XAFhbeNztJQXGWhgGk94FIHksYZg8tHJaDzwblQvjqTgDsVRQfggR9
4ovD7F37ZeHpkXSARFyLiuvouSv/JmJFbDzkxdDw9GndS/4ymGH3lirVzf3QgLbleCy8Hm35VRCK
QQuPw37F+87mm9Sfed3gb+CqqGbg0er0ZxudlvN9D0XyDjWuAx7N3B0Bl3l7PggtyAkEjZtoP4Ks
DcPYjrb5no0hEpSXWHI8DYEgSOLjnzv0y9dbE6ogkB74i0mQvq9GpBiOB3VvNuHmUFbF87f3Lpff
7pwZB7TTz7QTxCnKW4uHFf1rPA/gM4iTwJrzeM1iv6I/zWoVUcipnfxqczZXLwe4nMdwfVNqdsr3
kQXzp4El6vQZuzRk06+YbvABrXqHozZvuG+wF4/HzEtfYmzS16ybDOlCuUXlzkAqMDLJW5u4cYLR
zZDwnTDhDnkLigBUZsAf/vLkHu2DyMNnlVB0F12H3bxkFn10p7rUjhyzSTBbJsrJ15OWzOeBl1+a
vYu3Hf7HLhMGo7MoeLlAOTjVUvvHUZv+gqeMBv9LYlCpnEhAo9vkIMo0wq0T6XyNFGnLGzjUj58T
UztnusbCX9fxvJ1jwTufTjsWiQZCp9B6EEyTIl8vBicziwhi+99ELEU9iUg5xFbV+4c6wGtHoeqA
Jdkj6I2t+AnQJAqazZ4RysbqM8XCMkzXUuy/LREBTicPTVnbaNrVF7RoimvN5BK1iAfwgaWzgjHW
C0iyrgNEAFjhfkU2AnkPTtdyVaoLReRemz2MV+03O8RStWJDlVXpFJoFK7w+NxTNEkEodpaQjhID
HWB9FUUZQ5SaEkzmF4+Vp0B8mqV346MCjjxEjm6DSsag2g4Ylimck/IqIe7WCeGISDJ8qI3QGNyr
R1evJcZhweI+B49MzQ3QlSrgdk4oMQUldGuy41rojm+agNhjFfj/bYmAP45wivh0byPQAKCCHQT6
AojAuC9bDrG2AW5JKXqXS9boUZsKts+JtRWhuNyctJtkivhAQZhwS8bUcaGpAinSqlpKABqUlSrI
ikgVyiyUrceHsVze2cEvijTvR6xqIkSMrKUbSUpvndo6QYwdfXoEgjh1aew8olmuIwHc7mh/nzhw
v/g5W4ZXBfXry63n8gY6rz5rOsKKv83eAGiosLZ/HelchZgpzcTC/UfNSqOrKjO7/s4qWTQImZFs
zwBmuUJa9IVGAlSuiGCD3CMJWz1c2HQLn7h0C8FuK/nF0NqggyKkKV/Ko6TUm4QvuVeGMXrNTeq9
OAG82Ea0uK53HEg+cR+TGLYas2pRFYR8t3wIQjUNayAvZqfiKL10HKnrCzP4mA5Ho8ztvxXq8KmB
z/u8exFbrpszaho6hMYfA/jx+nr8tpys/F7f0GLbmZu8BR3LH1otv5d3TaFBZyvAh5+SyG1T/++z
ChvUp+yDlHRgwt31+qmu/KiPvTqV2vvsZUfoYGIzr1vCeg//0YxCFZaMH+ATgAcOWaehJWLDZoXk
S+u2MCK9ZPr3GrEsS1zNADg5gE+mJjgX7iG7/bAwSnXv4OX29xc/Rm1J/raZID++M1DAe7vy7g8t
WNqMSeloEoj4kcQHSGTu2OYkB1WHgruXw6g1IJ/6TKO7DECB/mrdmEQjGaUXr9+yKIsJaEeoVdyR
ZQXZOxiUePCLJWjoe5HvQS24TFPwk2e0jl5rmjNvOvkLiniIuLT7G1UNhWdRvDSfp/wkeKyOEK5I
JRKNfWDA/CVi5LSfgHMNRia5LX0kVbzOB3tEvgXqspjpSW2KQivV+ei4ZMVIOBajj/pJupjmTMzC
13Qlnc9W5rEc6HMMcxsiAdbVTTICYGwqV3Mfl5l1yzCIFGziRk3Iy9lYkhw1CJysPQlIcX+GxvI7
BHnga0dpuebTm+sT7dYMn86/9/beebMV1m1LS8vKe043gUlZ9FsbdXiZxKJwf4HlU1MzKPudfuvs
ygLUN/pJoCcD1HGFkZSFy7jj1qk4/u7Yup5VkpW+tmjJtkGDnr8+T7APHvNbgNFEgr4cY1pszWn+
lYbV6/W6IAwJOJMzGdZzlnRA5EA0HHoJXRzba/FMCVLsKfhWTI2fyHze/8OFDpl16gAW5pmP8tvG
QVStKK0eL+vyyxa722OfEp8VbTmBBh4gFeGAtDlwph2irt7X3Ua4nUmAXoQuUlRBoXL42Fya5yk2
CFdSO5rp1URmjUAMF5xXqxvdMsXAymZm6WqR2YhBFxyU3Un7qISBmLczpOhWIy85MuK4UL1ZQa3T
pLtBxKD/PCrVew5kQ1lWXQuSrC+Kh0C8qAgui4RSaa88I91GYiDY5WsQSHQqNfa9DB3Q7MR20z/5
PhTYcGYNAnIufYpHndLjD0GCR62au3e75vhJAmYBP1qyrAY5sqOyEZHkHM7WY4ZX2ZItQOWhbtzJ
fWs7CTyIqSunycwk+t+umkQoRYY7oL6zdP0ruYziYzSf71dmECU+/2MBZu1atvwN/rKGoARgbecA
kC1ofnO4IE0ZJbwlZdpeNdFhZ7/QYvgYGlfsfCX2vcJM0a94EZHFpl2jdi7gdzz5hfHr6mFabE6D
T0j6Jwh02i7CLdJ8VboCUYlNtXP9YWlzKio5xB4N2vVJeDUdEE5v3qxzQwQ331nrmNg4xB81SmlG
0F52JGPlyte9CJwK+Hr8T6iPaTA8OFiF68ngwu0gWgQJjjM2ysZ1uoNhJ/FDUypd4yHaWN29kZAA
tLHICWJSCFqRNaFJ1hx3hS0pec7DgoV4AkANBeE6S4zZkAseclcrtcHM4P3gR70Czb7HjcZNCRkz
L5yDFgpWOPTiVDOQJvv6jeZGhNvysk39jofVXpsPWVV9AjnA6EjK/FD3vrvFjfA4FJXuu2pqK3UH
v0A5MjwbhoW37YKpZ60bV6mP7Da+BuzU1/wJMZ72xAr7e1ISzfxbT+CKrWpikcgyEGFUDugmcsi1
Dc4XAdcdd9ABBTUuUFGtdmTVqXicMRZCZuJ+MspKZWlojRaGYj7CjfoXGRUjo1DAKVtMnuqfRWK2
FeBA0kBBokBlQ+mxy9mLG6qT1kg3qvpapFeRdHtZd6PQuTy3Yr19PgIfn0OAh70lvYrKfwDIt6Gb
xaHMTI4qbdlK8wdHUr5sxRwDlst1q+9qqwf74zkZuNISvbl2WKrRVtr+9U0uOATX8zQlN0kiVgQR
XNLeom5Pk+Jp59W0bkDTG5PitediCpO0RB7VGHdhRqIVYS/PmQm3q7ygFdC5JDcNhJMdbho0UBkp
BTgQgJcV18/HyvYmhiEEOAzvHKp7X+BMh66iXsw47nBe2B5gepnkPrW2U2mlsbSvIlQR9vtRZD2S
cpB4LNjTK8Iw2sY07/YNf73nF88SqILISNqiwmcdmEmf8P+tn0+Ytu7EmFEalzDnG0jLpZ4mq1mg
x5TlmcOqA/PnrJjnbpSmZrPS8B7+FujvrG+BDrpv+bdBCHch+EpICH3CAs3HsoAXuVEvxyGNfh8o
oxfH6N2sGRNFdLSTMZo07c86DqLLduiyTfsVv9V+bQur7hnuHMs9YQ2M48pWjheB2gRKVyHs+md7
PkxufC4I2dMhe7LhveV3/gFxDRMlS+XngBq6t3jc4N218ofcr/KMomiLcgvGcwDTQxE+fQWzRjhw
TM1LtrOqqPWPtXSKbUhzqII1vg+IilqLxgsJ7pdJMAdnCtzQcC2CVuZOym1UBgN9lFCu+VB24hue
TWDcGhJRC32DMzQnidmwpoEcMc9JIwYP49US3+x6TnMyzAlpq3myw4mWsK3uziYoEChHsNmWhLRv
sW1LEPRMK9E90ytFYRm9P60Ivdh6uk53/gB1/Lqlz8zGNPB9DtcXGsCBQj+wO7mElU9hIHoQ1Iz1
8fz/ZdLYuEz7TQC44qmYGeqnYJ5U/vygHWspNw7N3d0OoPd1yFqZQIwiwBc5mmdTSAuVHGnma5n6
vk7RCYcV0NuFuhu9PcY9uSZwlpN16ZkNXrMmhMtxNBZDxjO99cBlPoraAa/j47soErFGVV9PNhqc
9yPM7aTiKW8KS+3NF84g+/ES2+6ZIEOPWjzTc7Zwh5XwXZm/ynvFwASqiU4k53cigtarx4ICSLXH
Msp41Irv4Yu1RgUUHKRBQSvdAHHOg8N5BLZaGdjL97Fq1NI8gAG/P0AOy8oRWehKs0LcBPHcW0tM
IPObiQltzNCJApaB5pL/ByQaqaUnOS5VOrYSAsQ2+qrWxjdwjKGmpCWq5U2wAeOMNtaK3YkFmTWs
BC2kFkVD4jxFuiw8Xekw6o6ZcOIF4YaSKMbkBUp8j8HeiY56dqHS3xKBSqm0aPNg7lxtLMXpXl8f
GqJtljfZDdlo5qC3VA75axfQmhD3DkbI6xYZnqHXk/FYIxuzJ2OIX04Z+px3k9JW3xSP7xkaXkXm
tqKwPaIhj7hwp/E2vi3PiIWALYKix4qwtfzf9yfFD7FhebHYStQg1P765jOHGWIRER9Fw44KkMf+
kRjwF96hc+9odgZZbvBxuJIbhD8kOBE9Ou7R0fMQM6jDHiW2Uy/2/KLfYv5CBGkk196RJYyoVwuU
LsdeNBwfAFfgVC0xmMa1PidbiGO3S6oSHjafdLjecAFTB/Ctx/EDZM4WPJpGvHW8m8QvUOKFJagx
2YL+RIbZkY1EEWrXKWmxKMWJ5ewQXq7G9wPlGxmvjOIhIGMCo9tElt3B8cTF2y0NWlcaMJo5wltr
97zKHhVxMP1N+5zaDuuR8v/Kt0lzxWFcSRQiUEATn5u4YNcqHUsaB7r1arbOFbVmL1uNT6mg7rwi
i4KNYvXNdGE13yWP6vQlVxYdte3nC6Qe1IxgIeIKxEWtJ27GT+MqsYCf3m4TvexOX54TECzBMz6q
Ng0eqBXlBnD3TIMKa7f6m5j7GlLhMJfisavtE9vtBes6qaI9XnF+ZIdzXnyX3d78mlZ8JLr7RjKm
TJpSg2YwcBOTSF+HRC4hKLdF8Q6PUx+G7JBj0Ow/3nw+Vr+mXKhwiu/HT7mDVpFHeQkU8uCEcv07
i5scLfXlu8tdS+36JsC12twzaSV765F4P7xfLSgmyugIChs6fKllfpw8nKvrz5hn3P47XIhorCwU
/nH+DittW0l+vi92zwuzxMDT8suiXjRR6vc/aCY0EDxDcZ5D+lE9W5nW4dZcxGqk03StDN9QzwXh
02hDX6dMVANttgz7GWweLXIJYN0rH92cKU6hVvFw7atI2nhkDFoc1dWlOKRkyakIME1pNjgExS5J
3XtDGhvrNZC2An/sfF7RdCYciK0fflEnq2KsVS03++7TLvAP7zHOb30BZDvTZj/5P/OtQdEDFUzl
lb51mEgIA33uZrGu8n2/ZRlKtZOSIOjsxPiBZ0x0LzM8dIztcWn4kGABzvU0rbUgwxpGxVxDdPGU
4cBaLbFdQfUuYwSAlmObzWcWeeoshz9XdcT6qe7ELKu5H+VLAull7bWIcGsdYAFYhOyNbqDVEIVj
xj2p7jfxkOa+sd1ZskOeop/6ul54B6aOWpdATn4r1fdIc7TS/n6NAGixSMP4gpDdamyR2cwAN8yS
wM9Gs8L1cSZsvr7LFkRgGj5bVGrFy06CZDGcPpK0KH9K5q5eMoEkJlO2DQn5xZjoNEOMwBlTrabG
ATr43napfvEEhRwboev8ITHwoAY7c2H+hWoNmog+JTxDjV7KrsD+W+9Kp703I0FbS8EWmb8iu+Is
tiFF+Ztqxl6M8tw7OUh1j63bs1HQW/K0nqDX7SHzGtNe8rUia1Zu4bNqqsfk+xRzhvAPrMxYNFxa
yC4PNtapSHVI21cTVscbUD3bxOZ2OkkU9CQIojaNGh0Mz7LJ77YIHxFMZr1AM25vd52p2fra+ikp
hZBqblTUWdbYqeVwUCNFa3obcvzi7eMPWdjzjeln+gVXZu9VZzqqyC5cAhtpfJsSVJ1+xvx2GBf4
WYzJ/tjvmiph5c/X2u9RpWCUvhWq7efPK3z/pNDjahUd6cn4iVYey9glwW3XhGB+uFHkzCJeHwcr
RllG1bK1y/Z0XrimV2bQAYjTNd4tBDWzFUyzMcJ74ao9ffpYD5CLRaOMEfaf6GtqA3oFuO/yynbF
MqGkavsDMZyGWJywZCyXCg3U696bJjdXDRoA0HB2E/ep9QnS8CRfo8Uiu4BHKweduj5gPaCzKeuF
eqHhrRXFLqZws2Q0M6fowoFG1bT6tQ6tGA7PC3Mw+MvuOBfEdHVa1SbWC9MKsyIhmlbxgG1IpC9d
lmUEixeCerP9pdSP9IkvHZyJzFc5d2T5GTmnPRDnb2+RZzUYgC9aIVUuNwNgB2PkxIPTtve6inWy
gSJQXnPXbVjtNfxvSF5Wdtjku055T39Y0eHC9xFqO7u9xtKPYfzc1mrpbrNZtp9UkNrxO5uAGGM/
sv9vdrkc9ARuxZ9sSsJRN4FeoQ55RbhnN4h365W2ZmRGyJxUExheGPSSZTNk3vskyfQfAL190S0x
loQ224CiVuJnLRmmjm3ia358zAv0kD1+9OWs5O9CkOQcmIfTUyYFN7BB0VMXvK5ZenjIV3Yuyd5S
jHyOLEyHdCXfrYMiW3htoQhwvTorO184q0+7fpTevggLDFsU+RIbbl1Libpi+lxVzvF8kgZ0iWh9
LmKqyufaNyQRVWfMnmfORVMnSS+DZxoSwIRfL+LPUU3b3d4kiblmQdX3FYXASDNT3IFJOc4xi8vy
kTbiyIV3FIn16zGHITa7/yioGsfo4tmkNvtJ4isLUcl1k5Vx0fEudSr5rCMqBldxILoXHtXUsGCt
ztqboA6usNEE3LQybQgYb7EglknpsJ7BnH0x7y0NUUZ6Ow77V9YUmlQlGwQNnjdY+dxOi63j5+7Q
JQ5DYn7LunjH6GUntsmJ+cekLDvi0s4+9Z+nrCHst6O+B1H78J8dXU+HXUmPMfcCynr9IzFElwu0
6XZvUAwPFg58PTwDDdx/Zj4/Oayjivpwe/pgpgjqs6xUZJjBgx0AbgKZxI8/4dXdiUcUoS7hXX7b
mGetsYK9/34NegO05bZ9BZBxRFY312xaRwemI0GcLRg2zzbWM3zouDNRVHOz4vkS2icy4T9m7EYy
4yKDThR0z7+H8YXMGLoih9Y69tft+IoD0n2QCuI+KpQWGjEM9HwzdT1J2Cdx8pAzWu5Bs+KiqC1W
gaIzim5L5P2cabA3+3jAqbYPfuXIJfi98JgyCCn7m/lJ4T/y004yfLdhO/tOoLct9RM7xTCtSnay
6SRnMlImpysjoZNjwrAgT4A0BZt0i14m1tVGU4qplOHIfptVt4iAMa4BH+txC8oo2WNIKwoOKUMg
7XUK/NEJ8uMJcIAvecI65SPQq3Y8ACbkvq2sfIuOu+1eyABfBelD3Vl2g8RfMfvlyhh5nnl1VMbG
vZ49JKdyQ32jbKfywl7wR8Ae/lCZTdPnP6khcn6TPO9fgmWYP2qUq6R2uSy0mvDS5ERcYhi1LPf7
WD80LkeGNng3P/aavX0mEte1cL70x/LM5oB7fWMuk2kK0O14OK+RI68cP+pTlIgvN04j9GiIXI1w
Wi7A4VQsAUofipzunB4Ee0YmEu9ARi2D8jdXx9OcRTb500xq/I83NNR5n51qeqpZdl6EjQv7+39E
bkzHaXoBZsZa5rR857bG1O6eaEcWxM77QPEO9mIcYcHTFRCJt6d0H/JgqoMiO7t1snDmQb08d0LP
Vd13X9GdDfn90GVktPu08ZWyFwAkYArHCCAV5+HpvDik5tRvHsyI4BJeLOaSIfU4WqoB9qOngSEC
4PiZbyytpKlH9T4r9G09aX7YItpqnThg+LqyC8s3Rcl3h8rVhcI5piqp4ANtO6LCAkC6OTFPBRCo
BFrpMcYaia0xH0MfvnpZG1fXrxproUUL2uoS4mmMfTzLt6QwzDCsughXV48Lyh+1KHi335ya524r
u6QCXDNu7upxEh3iOqeArKr1myVm8zp81LhYXq5mVezqCJQMHY2iFVIn3BahbVBarLgjvVNo3fmu
LnXjIi+Bk1C7tR7fDxfE72i9JoSV2517qSJ22qjRawvPt0Q0Txv3GmtsCgZoSmCWETqVomiYnkQi
HM25q6XcRQuE4un9cRqco+XV6O8akzflGXonUTMaLUFfziJWDOvQrv/SzrjxdEevFFzvMou9+FEK
zJNYaOhTzKnZ13LxEfFUqPqQr8MElEDC8DOsp7tQ740gM52fO3WPE84tP4G5xsRurNkOPfBkpk4U
OvGq3anM0Vxnp4InD2deF3Z9KhUJmnXhX8pKlcEqq7gAvQgzbM6I4uI7jEKEhwhtjsEtcPKE/PzD
y3eNOe2wLRTNQeVU13B7gGtJ9hBcx61Ae1KhquFGZyAbh8+upqa6rqxGH2X0ddTOEyIBI03mkGns
fVZ26OlO8ABYW6ulNz4oWWmuyqU+MQ82NqliQmwVw0q+nWj+/QQgDu9xWo/XToisUy0I2Skb77iH
067a+xe3XV3I82jl4NkUqDwlLI8nvn2r2D2lt25YjHNG+qzyGwojB9XLKDk0awZs/d7AyFVhLF9t
+YeFRdse1vIfLMoLD/5KrS2d+WlI3EDa8H+hFHb6+pb9TIOMit/Qox796tt5v4fGa2neuUL5miNt
yHd0JBRDwGhiV/xWbbSCJXhrI89UYoV+Gq8WpPU7XT7NNHSUzq5RmDJiQsPekQFH5gP9r44t3qVA
T+d3KUYxRHolwyV2idOtuuxgZRyj9crjUEcdLP3NqbjYuHKz3azdZrcNgxmZuucWHpPMZ0sKcRTd
xBrR/99lhMbRldYipK3LfFAAg2xiJDu/400bJXsYm/ZhKEBBpo5XppsojRqiGndwhV69wnCmOC3e
vea147/37763tU3CwNz/Zm/aSOJKQUtLsHB182wpOxd8YEvsVPz8KZlSi0h2vHtvXiJaPBT8+Qip
xB0LiUjSbJHdDXlSRUC1cFH9VfWiIWcy5Dm4EfjLL4DmO1vBZJ27tuPWtdZogYQrB08TzpcM/mqO
WDwMeCk5DDVrni2Z749ouCMy57x52NINX5T14trTyGLK/mS9ZAziKzBHDfvBap++HzBosuvGaYMK
bgb/k9irEQWqyHWNWH+VVPuSy00B9PhNhELJz7NCofijs9/9qdVCzFwKATn/GqPnqMGUbek5qCTb
nUH+KXwDz1dybrIDgjuxXYTKYpqOwG4a54Acm6meaomVOMvdZdIEMK3uLWjKHjnolm/3fWgmS5nQ
jAtP6vE2MeSdikCyvPNT0++A0WUWW4vW8zpF3jPOjyv7uQgp+aYZtO2I49dboHFZfyuB4XE/1a6f
tIdIHsIvla9M8wH8t2qy0eop83MCovPtSquT2qGZl5oN82/Df/6mJPmb44l429jXE/bCOkkwB5Xg
jOj2xWokudvyHVG/AKEu05VmIKOnOoiTtgEQDKJTLyw/IxPDj7kBQSRj0JKQPqd8NL6vSII0kk+j
TZ6JExNYC+Sx8FUTrBG8BZVDrJoRVleMyPTJKC8St0FENeqAvjx+pfcSI6xMIyDip771M5feDlIT
8NkwK8OeJ3298uzwg9ZLuedxoK7jXQ5OyzSqyzVeihwiU6BckyJ0UfXWVn34j9NGd2N4XgppNEP2
wfFP9kcLYQYCGf5MylCwlEViA/IosjkCrYuOEOBboeE73AZOdjKS/AEd3KiIFt3/qUYAFs9qJGHE
PGYnuCWKgvGwUTpes9MvG9gpGg8VT6kgDFM9zXG4UwiH1apNPUfQxp6q4p7cKrWRooSzYQJzrh6f
QJ6iv3FoFhvHIzU+kyuZPoMBSarSxWdr4xGPGA4nrTWcNMPUvgDG3BEv5CUuAfEeFn+XfEGXPsxr
EgHFXXhydO2ErvFSxnj8FEsVQtcW0K06xhuGbll02wJxp4MMYYc0I2PDWSp0EQJxdH9G3BGWi98r
R25hUhrrQf6tGmDqnZSC+MbEXP5Huvub1eJzyhH1RjLxTXYKimmW5MI4NKimuDDFvRP641Nz8b2r
niWcmOo7ZnNaEiDbMZIu2pURX4lYufogcvpvKnKLJZ1Ty265WVix8sJt+w/lv4OPJHm4yr8u9ZAu
NCFsyPflknnGQhuAlEkCMonjVB+UBoHAerQ0zPKpxtfaFTwAi+hjtmmZLA34LtveDSzJhzEw9xDo
LgI/jdCFkUcOjWddCcKIENnzl6bjTlF+YDIX8g/Jrf3IDVYBf2qPsuvxirp2L8MkZHCR1IvKSHfZ
OTEOmoepVEFPSYow5e/16L4BrTKxzlg4v1yopD20p0LiUbOTr15RxEzqm2N9xPQOAMcY965VbETk
GbfwBdVKnY7O7uwiqAGWxAucwCDbF8/dda/sNmPXCrv/JFm5faMi+LQzSMo6Tv0wnZpHLhHRjCEC
MaxN/WLMHtYvVqFoxw6Hrz9+uVmB86WuZWhEhKpmKA4k63kh/pJw0kQLdv8dIY50WVEbL3+g347k
JnYLA3lh14twj5C43f6R/kQflnAiKpOwp9mM0Heysuf9/TXRyMRybXK/wcJqcM7LnPNHWZZWYry0
arFIectDeV8dBGYEBFwFP/l4/QF+3GMjGxgq5k//vHdm9/He5DGrGP5+QUJrTgxC9hVuzYWMHzd1
6vDwTgk8R8PkPiITzUzmiT1nXFDVymWFJ34VyP82EjgTq0cNPBza+Gq3CBNUKIbzqqHwcZW0WJRG
Ea2114Zpis3QLwGsR5+Ey4nFtNg02AXGSmx+nvSkgcYGjweAj04QFPk2EsTSInN7QyH1vUEsVQ/Y
cxZhdxlOdbCBwzTHoAPsW2argOl+AuLOWJ8zZGBfDm2SVdku69pKa/jd2KW9uSzaYVm0E3toTquR
4ht2F6cuAaZtrfdxk/6UA1xgIJZh4sa9IkgxPkgvPmIFyzXWtC9EGPBsOUlLtdOq6tT5peTFhydZ
+JrvcQyRM5q3Gl+kk0lS75Mb1HfXG0huxKC1qN1R2ZIw3mMt8tUDlGGCPpfQE1kD2XnpOPsOhB0G
TYkfjZDtka9gueH0Mm80/CDGlbE0VOQYqSwOJGIQFww5A2lypeVIEqAD1KP8rMyEWSRoY6gh7VOZ
6Kf/4zM254ijl1MnZiJJwdaeywpmvkkYuFNStfvjuSoKHd5x1IH5dqKPGX7FmQsvU0sZq5KYcbqo
bhNL169VFZs/g3s9/bG/Ugwv/5a5CogmBshHtpi4lyYD964KY/5QufuubUcELzq5eZbFw7M2FeAa
9+OPUhlxtjABhRidWeNU3lnfiG11JZ8YzJgwIkHbLmotyuXP7XEDaJIjDg4pNgN4FFRyFTAaQvAw
Aon5FvBuW/wT5bvD7jYDZlbk8d1sheHx3Y5yOImNUvSd/sAym6+GuNIRQVD5C2lsKtIeAWh5Y0Gb
AtTzdjopgFUxvWvyDRCK5kQP3JaMFJMC8dOvbQRwsmb7ZpVbpTKZg1FmQN5dcaEjFyWoAvHM/BCX
UtjX49pHJkQZS/xH+Qt2wzPL+pLhfBp8VV8v78+rWbmpWaZZQp45L0a4ipnTmVK0K/1NrovMk5I1
Hno4HuSdHOZYgjnvLxfwuF0tWzego+1cQIiugE0HRQNDzlaoce0iDuffhD1Cy6P6EEse8Yluqihk
A4mfQeVvtxyMs07S13Jis7VcL2fvlfEqnrjyYHXIwhbKJmerPAl0So5CzEZGdyEqRmcomnzJHKCx
U4zKeTX9BIkDkUhw7kGVQtDOr/GFpXXYrlW8hYU4VVPK3OztW3RcFpGS6WNiMzXO6xwPvmyzIitm
M681dEqVWzynZTxlX5/7t7MsjKmC/WCdkOI6aAIkecqIAmnTASO9sXLBkbVsTg+qzr3w2RBe54CH
AQmgDqxUcDQpU5/fmVu1HPs4EuSb4gJnTsRka71xJfp2dCwwewaoRt983SUViguHAjl08n2toKTD
OY4ebGnzs9q73Z6ux93Y37V0dH+ucC+MR5iYwkNpRFJvSpduQ5yz9XAc7Zb085z/k1WkSfEjpLpB
Sy5EPdX4FLAos5hTBe+RmWN541v2YhSfrjdHFevPCG3dJ30p8NbNli72yTfK7ezh3BHwY4+px3II
H2qyGY9bpRMZdigX9AFTD2sHOxElYpE/Zdmdr3p0+NFM+vwR5bq+Qds5txUQBQjSi+MsZI+bxXdJ
7sdDXc3i9LNtum/j9GN8VtG7xOdUBOg7auBAeWbBwx01PVLMZBj4l3ZTerXWvq+opX+0OfwlHvEY
CxFjZ2XqMJyyjk0/GPIi5YhHSXtDHRarHn0YtGEh30x+/nbTi6w5PWacZEg3Qyb4EZKrU6pEe4z3
d/vKJyY+TdjWAntcGHiIi3znMCx3w0CyxGWOCjigw9yypQVaGIoKnE5W2+1QcGFP8te15YNqUqZM
MZUNMpmbM3bnbgaFteNHFdjSO2/4MN/Cqe6MyeWhEhyD/YfA2mDvlFZDS2A48jETpizsIssUAYIW
hBY8CqGnB6z3nHgdLLpdAd81CreFih7Etkls/dnMWMI9FYUx+jqXD7Xt2fzDEcmXJIDsJpCha30k
ZOdx/kihTS6KsoPUEwtQxjtngneNanHZ2D+B6iulWqrezgYztTH16Z/9qNb4WNaB3ReQ3VXHJvp8
vA2ZH3rFLxA5OCPBJwpcTMcKBGBYKSMneDylJIx2nuBiOxZWSeAj3tbwlgQ4rpUiyrUhRzGgpOmZ
CWbJFAme+Diz0QkFpW8VKnhjzv+Wxx7+Cn3tuLrN/oL/lunbJQ4wn3XmiMXARLoH7vBHBH1WvZ2r
II+GNd1FibLpf00J5H5uIXymTcF+tryQzIWsWL+a8ervVkRdrSvkfh/mk+bG4yCMCU1VTsFfwbYj
zEimeLDVyyCuR80v5QssCv9Pkqzn7B9EIPzWJMlA3hqgL6Ji9ltww2eg+GfYvmmOWySouikMJyuG
CzYlU4aP4oVbs8PpWr9pNCuVQFH5+E/S5cze1rvUnXqHbty/xTOyGLM9gFIv4E56gv1qZA8fRiWA
IV1+9qD7QoKwm0VmqpOQXeyCM0tM6odjkqyaS+UQmKdEdf4nSxu2Q07v2Cx9OCDn/vOc2rPHP5Y8
P7I+YA1dhULgLVWvaMuKcxD3ci4VhAUnHX0PDKUATNH51O1LeUyM2IWeOan61qsmhYiWYFdRT0La
BVcQ1QdCcNdA5zF7E5u/z4QLgLBnVk/pN1rDRXeL9fKUPhbd7n5uOvX3cDCcOMgoFgy2qMuskhIQ
6XeHAgA69QGHg6sKR0bcbo43shomQl7V7nbUZzJyJsjBkPXbGgVyVXGP1Cb/XdBXgIuHrkqMfBHK
QuLkGzDXKMiCoSP+Y0wBhdvaaqodpwxpKc8AgXHUUI+HG2FltR6enOnKTmYASc+I0ya1lsc4/21u
OSa3XTSJzP59A7AVuDar+SOQxEiedMeA1irBXT0aNsKxOKaWW1MyD2ek13bWagvc2ljxXD3uJAiy
7Ra/+foopU5OHXzB6PCPob4sM7HuVtbgc7dO4SaeZFtjWYT9U4Kb6Of4pveifMyBQvw9wsctjjr9
InI9LPZrdwaVBlxbnwecoruXXj7jKRkgS1xW7BDr6Uqjg6wdnlnHe49DkqavJIk8AjmEbz4W0Z3o
SZOI5lxIEMGw1PHZbjxlAfwl6yOPy4z9VENZ+0TPtitJMsBrAM5Vk9/6o54qAZlopfmSd13OBQAx
MLUyKOdRMjM0yRqiijy3cSTaDFJw+4BNxik9AOWmnnfSN/KkWnvU1phMFHizMMTHYZdNqdLVrcyu
8/fNpiIVmXzMMUmzYk8pLkJnTzWnN+9ApqCUuIC1ZVpSCyMWi1JKAuBpewlhZViZccTiLiEoYdLE
6UcbEgmfrm9b9eJ2T/2ut29iKUMI+vD0/JEXDGfJIPE62nDe8NZzQf9fvU3WZtWGe7ts3FGynvEO
4NQpzaYa5yi7+rZvQwyNrUD5w/28r1F/VIdsmHBQ+OLvGxL9Y8ZIkBjt61q5WR4ZbXRSE/KqGYCO
zfAakt8AI5osDzn/DIBwyn1l4CKDV1VcvPajac85xlB1/c5GKlV+YfVewwGRts2ByCKRSQOA+tyZ
sFcLJBL9CT+aZM/hqNnijQhgyXxwRCqhUM5Skz9pQcRyK7iaT9cvXfU4whi9Qsk9SQk3O79b+aLq
IzBrJj88yLbxv1xP94HoJqYwhylIHJ/g34cGuYnH40cIVdXoZjtNTJbsjM5H9ClrxHeg0DeESaiJ
XCudFPLJhCbEkYcFKqRznTalD1aUGe92Xx0FDOwqwjUlVMjL/ySsX0B19cRI/YQJf2NUX9VvA/+/
rpFMPhM7fGHQnl8jbMIfdEWisyQVrD7rGgLKsRB6/Od2UZcF2PrDS041/qMBXRY4QZJ3gYPJHq23
8Ss50+rIVS0uUwDEOD6kudyKs7tuL5YG3jOi1cpxX4j/Z26O5oWiuzUMzX3313AXt4SnQgX0p9J9
I6nzXytS48Eo8DDw/bP2LQChgVEdgQBFOCiIA3GtF9z0utm/ATfHVKX99a0BCB85/zaiwk72AW7F
94JAmCZo2SwyxC7JBLZVkE3qelN6hmg8pwnT2eMkC+hJAlEj10KrTYBraUA4rdkIpk2FjRmr63zP
AANexUMMRkGZqwVz030A9LBh9OBtjz1tjq/6TCAedkQHxR2dvTMA269fUF6ZGdRrzI+yvbdo/XFA
4SVBojJEjTi3zBn07kUhjceyNu+yR0CDQeAnq10bcP58tj+cE4NrQohQJePBsx1WVTxqf8iq71Yu
W6BnsiBIt/cdnHoKECPzOokrMLBttDeHOAJOyoAbQncnbC8DNloH13wW3XoPAW3PUDUU4ke583LI
XhDsQyM448uVZSe6V9M/hobBaBEfPEbITDAiAyr6V3E0iE+1Q0cWWZ5QdHFxv2mGyj6alrrfiT1Z
JmMUYlNP95tIkmJY8YO9xjXhSyXoneOL5wLxQVbNcYuz4nRvvWO9au8N1LmE1kpFicK3P3F5cN8T
gJFTzSY2ttNS3sMULn1KNtXMo6g/Tez+0LE0vZXyG/kkN4Yv/2jhqzIszuwhWXWq4H0F+H61vr2G
7qgyRmVLmHeMKaMjftj+HT1opf/7iE1TyMShUB1nRUi60dZMZc8jrzq25xmvN7kHrrz1pKL4bsX5
zF82c/ns/DUB8rwHKq9Zo5qTI+Vpe4OmA2u3eF5kPsg3QbOhGqZAk2bf1Echh9/SxGYbFG6URJNX
ExUyf8olzUDtmmsdohdoB0jY7KZ0zWpobAcoqI5pDhM6PmV12PtlbzXTSmCWcNQCXrEW/ao3JwGV
UWXvmjZMLvbvNfmYAM1UAiv4aDCjMshWpE26TB1UBE3Hqp5Tzqm7CzNSJv5DGe/ZmN2vUEPbCVvv
mCn1sVC7/du+0uZYs4J/oNoN8d501gOE27TSkQM70+CWoze7p7nDgraIvwrW82fJulk4ZXgp7i3K
QGXivlbOT41wG0FBo2VW0lLL18HyzS7UOnqzD1/8cIjDVZNsqTGtDUWTPAg9cgw+jwjgpCMCPHZg
vtJxT65h7QuEaIjwsCO4HxX/MbWRZXUohDCtQmxljlql2GFjLWXhh7f8VS8IFGUY2nn0w5rr1Hw2
elqspZHsqy1XgFvVv1n5x0c0ST7OmiCngShItsVUBb3leMCjtuSWLeNnXEnbGpsZhrvcVKraDvtk
SnQGKBJMtWpvltP92CgfwvGw4+qOUQZOppRWhyL1UBWmMjhcfcSTpc3/g93+hP0ud+o4eHVlV/dl
nnnOM8fvMJfdcsqDzu4dovWSOd4Ab/YRHJj/0O9BUzdvXqdUpFgeGslbWVmYcKfe39PjBZK0BB70
KCj3TYdjpIVNmr4F21vO+VNBD1gnKKgdzV9XOtxjrP5hkdEhd9zLqnRMXrfSquYNqgrDFLiz72Xx
Fl4wuY9eQspv1yJXRdJTY9rR5BiRn1bDyw4/zI7UYjWAS6Nk5uit7Xc2jrC+YVculaAtzAZk2LZr
35aLmewbToHBmTwBX2kMQJ2pVQsx3yPYnM3HbD8XQn3OqW+u3yrC8zeLAta09JasLG/Tz8Z7rs1G
h6jAD8tgY2aWJKBu6A0yFENEKrY+ovLV+NXtUndw61kWgyEemUeWWQENo61ywmEivC6C6EiOoTYU
cPRlF44wwNQavL67VYxrXgdIm+YjMjo92t1UJJimidfz1GrvO5VXibdVvnN1xeYaKdPGEtDYvNh9
RQnZQwFWvILPbuojOFBKKfrYNKwnhzjVPSAL9w4kHuGLZQN5jIVjqMc8Mi//QLC8lS2Rpr0wVYME
rj+vrFQjl2xCNmj7DBEg4MIOpRM7VvIuQgjLEVfMIO0IaA0Xipc2AzeAr1vRgIV4Yqhhxt78cKu1
FklR43b2Zs468NK1ENLH9rvaSNfhA/uQ9BicZoEXS8ozPMq/QZ8LTqe6/tPYEZ6BiX/I0lgfLPqw
BtJjutO4HXda7Nm5mCj4VLIhYSSam5UEP+gxcCLnTzEBkqL6La4LQ/IUy/qWPMMa2+Rc8CJtoMNl
NMmkjc3+mRKwQJc350nrIVUwhjKY8t0TowSROCbGXKyGTGtKmYlMfCe4UBG283zDBuSMFHi5I190
KsfH2UErpQDFIqSpvMX3CYYN/FZYcppEqUrLKpUyLk3mFMZrjZwiae7DwjXXVctOVISpi7hCfhkz
vt0uhXmWxkFmnJuVo9fggu24WGH+gf2vx2deaHc9WseVKN9XgmqsZbMVB0SPXgal1utsgGFMstv7
Ie5YEcjkUSj8S8+PUAlkmr0Go92LUv3nd1auHIv3X0is0FOAeiDMtcmlWtdsVo1chKQJorQS8YC6
TshgN4W/NyRbpNcbAO+W1khALa0R+FvPZBgctoBBgSqe/Laoe7i8ndfggP7w3OYElO4ILbOOHh8v
u4LR9CELobdj1fVPxV/jq1FJATHrO2GtZSByXTRD89+3nDmBqmolAFNEP6FUk5vg5dVJbkizVGjg
kHBBBe03fZtd3/RA7znhHAmsrtA9yV8WQDUqTgTmzXqF6QbrNc04u8pdeQ4cEeKa3wh3PgSS1ZTG
AbW63fhDW/+ZXZBJ0Y9m4haur8G//UKZfN17H9gpOSUwvfyMy3odovtUowwa7T32Hybqarhp1rAU
UMWSKW1Eq/52+z/U7/iN20DzoZOBHu3nBRmv47XHYC3b/jaAGf/Mep7WefqQTdhZ8q5aQokP75Wt
ognIvRkR5QOxjJyAql2rFRqWAjLG9p6yUGPAEtO9f8dz9GQ1mU41W7QA2Pm9avHIXKce/GnfCHuO
5ln/HhhCjDUVAbE0r2yvKgVZPl4MRs9apJnPHesqHyhK+GuW/5kGyqQr/noJMqzNaaccMLKHMY74
oCrG6e4ZabhAxIhHR8vDc9ARislFe3GmDBeJBW9WqZ348QrngntbPiAof2N7CDlHcErY1bR/zVmN
RkrDMwpZA8jmB+A8HUdyB/biI76quj1/mPxUqH1T1SQaKy8wNasjSHfTrb8dr4NT4DCUi8Dxch/D
XVvAxTyvdegzk/YZJMU6MvubEGNcKNAg5xja8icZzQa2ixFJB+4OUPNuk2PnrKFIFj4JxANE1BTZ
KnT0mKN2oKpgy+zZU8f8NnpMehpWUJFmbolm9nfyLgcRNdg8xtpw5OYPyPAdKXq8qhnYEpusQdjE
LhjMDGs8O6Y0RPdLBtTH6ddwDBTF53Ik8DRzYHU6116D2M2tvA9Z/wl9QU0sJ+eV8KMXrse/LMWG
OxjLy7eGGoqEpSkLX1abRvVu6xvF+0DRkNWHk5RhdMNrPnqUEjEdv+PYnkisz2LqCTkzFyONui04
VYsMSiiZKV2LtDoCU9WLNCmDQEZh91SrOGmFBbk7co7F8n+k6nKnDwmnqJs/wYjALp5nf50ogbze
ui23NCY9xJYH3RGoDTsXH2Y1J5BGOun7ENx0YOqHqU599acijjs76wqcfVlWgOTMFlpPLZCL+hT9
xOuSVd9JDB+Pm7D3P/GHZ8s0Qwka5LeBTr3Nqsh90tSCY1idcLJhKjTinP1qU48R/s2FgGP+y1ci
UMJaHuyp+wQHxYO1xNaRf8698vVCMW7pVr9hswmH8Vnu/Sn6mq+O9qlwUDKwX4sQcgCT+nGn8F2y
48EOhGLSGRB0kMllJn7QXyJlvjdbZzVOuLpRqS1fXYzRgxqiD4NKjKTMEz/A1KsKq+p7RfFQYgX3
ggtFWp0ZykqwlOirZXHbpKoBTk9OzjwY5eQ7wTkvY3+2QbRjtP/seNLVCmw480J6HWjziA9dnRyy
xQQ/Nm2YR8KL/augeLpwRgNcrZ9IQsTY6ixTfBbYy2GZ6hhZdY0FnL4gk4RlOJ4Dvfdc6bIcnV2w
63wPa2UffSMCjKtl1pU8IVXkvJK3080WHkad7tBSkXPoHzxEQpPJbFy3eNOfK9+UnULoK8WGALN7
RSHAic2MmBPgvSvDlPDq9d9RvzDRwejZlvsjx/kr3eYeXQ4hMgiAP056wUNMWcbvkbgHA88qiOMw
SxQBjUfMQY6lW+gEMRsYLdrZJa1+DKnNMJ1eT6KVVy89UoREb3K6rynsRfocifeZ+xy7/LTs2A6h
Gws5sW/co7hdrP/9DDcjhQSpSvHfSFkmvzj+ueIbaTK9INnx5dzd416InQ9LfNErY1XjdxJnd7/o
3reORUt+jeud++NvtbnbzArUDUMPPssX+p6s4odnCc3i6azcrlqLd0uDPn29/lTUYUDs+4tOK+TY
N8aDC4Gp+D25BTGwPsYwVudqb6FdGxK65xmA1LcpsXquM9dVWYFaugSz0/6ur8DE+8xgIQQ47Cou
4rb2C10nkKyF/BBGZbtZOnJ9HNVHru7DNwGk4jgxjZAyKIg25cXf30kxpHfv8gkA+aqtGgLWid0R
66fHZVqCM4W+JpgmX84iVvdlEDiQXxPH2CITawoz6E14vW8B8uTFltM4tkR2OsvjWLay9YtULnzg
9yD+o/Zt7i+004SR8heABlN99HnQ8YYyla4cvIEIrPgawHdZ1x/6CFFuuZWKCrqKmyDwZprX3WE3
Bu5v+Ga5OtxoVm6WHMJcFE0gxGxgZGSzUILpgUpPubcEydvMFMEzBGUUiqpgPMTUDp9aPZmXRnse
LkIxK9mkbmS5vwX9FnGUjm9B/wafUS9xplvIcF+m13dGDl7dCuQVswNi5sDWllUtNEwJrneyY5ho
27E8LFMO7F6xjgITo9iYf/1NKaanNluMgEYLC6P2PGj+jgxpEyCSStCMAUOL7aG8K1uZlcBhfij5
3CDSUIPlfb7zoqGraONVvyktzwALfgBOOf8szg22PhtwmWfRixXWgaFGudr7eaOEkLivoP8PbnfI
jXSu3MiFFDfOO92KnyaHVTrv5C4gsKadHTFE6+Vz7qcIY9d6DK4wYwO1xZ6LAQ7f1pqDMMntZyvk
m9AY1M1bns6WpBCZNTRLG1rwbnC96ZV0wlbb0IXIJZKa+K0THf649BxzRn8QCCOORiA6kvZk9NI+
XkPMdr0FObA98sGKozANi/EoyvAX5qvvktb7wmX1Apz32MLe52ZTd5AVoeeCeDLNfFzOcfsr/kdb
X+LHwqNHnpYcoakLedHMv4AWAOJZ7J4TjWgNpUj+HlskETu8jvwalLbwSusdCLtkgIlboAw7/0pF
WLaI9Z6+a2Js7aynOPEXhAshZQ9XWZ9FWd3Ln39nmFvwkB9yEUHtvgFwUYb6+PDjQfR6EIi0d5c6
Wi0mzzvw0WCfzQkHvvVNmIpkxxrrHM+rVCMW4PhtoX3P1QGRIIKv7nHDjwTGcUewg9dAWJBZ+8zO
YUmbAgTQQbnNLFcuObrZwIqhZKtRPiscUY5eYFxLGVMnccoay+nL5cXlARscMi/D/4kfzhDEp+rr
PUPaef4SHaAJwB1ohHwSsvprIJTjoOi15J6Abaz+eaUROu1mXAJuSZQkbUjt1q0Dg1rGfh/Cee86
w3rmY2d9oTqg/aY+0cckCKSjxnK9Vveuh1gnawym81sFBryIQGQnJfKKrRuJlRREd0y76kUzhoJe
jWEpU5AK1ArXRjjd0ZDGY+cLnabGAZBfE9cSa1B5bvmz6TAJjQ3xtKxpNR8BXEUJ3yt11vOWZsbn
31nQLuBUHs2hrmER5UuMkYqDwkYLf4RXeir3kmCziOe6xmVsSLNjlP7O3GHAdzuZQ39gqPtvg2sC
oQPmo00uwia71CvFis04znTsfCt6beBgx/OuLS2m6JNAnLZg5rD8T5fi5J9kmymigT/j1Mxj9yvr
RmJ6gDy30Rq1j8vPHJ1LTdMBF/xVCV//LFSTsHtw4Co6Q+fiznZEXbkX/TxABx9BfvXFBZJzfWML
SacqXKZgVMRCia5eP0AagX+N+ZjYIB/wXxVFKdB3QJfr1WSPMaavCqZ4/AKHsDV7uCh+Cmdz/9Qg
7vODDATpWYmonyWIpOFVYHnxcOCc3kJCuA3Z/479uG29kppdRvr9NYzU7uUrF05eMZA5kl3gzVgP
FK3DsXNQwTywi/L5QV9KPmcv1Couns8xFaNBu/BO+Eq1Q813XqAQ4piwle1SA3GLN0wPl0qyrpch
87s5bm8LHdnYKj7HEmzi2MauE8r+D1cE+8pB1W4oHPm6zq3soBFy/86/+j/77ajVCp1jGvWwfVZX
nzedZ63wv2bFpAEnwy5eIOjZzptixDWWlMb2TcWD4LK4X/8nKhwUGDJ22XD1LhdTIOWGIO4qEK63
qBMfjIEtPod3AfH/vM2by4OhVUQ2/eiot1/VfZxZ4s2LKpWEsXw1i811JO4PNbRnNRCFfrJlA0Dn
0Olp+omvb3cTjKlfJ0LmWFrSLeYt6WwXo1iuqskBc64h2B4iTWpGvQfA07u0A7lyD6URBVFCPtbR
aWg1e9/YXCr/YP1a2nPLQspRPQmDpX1aWWu6Xx+O1sNtZdUBCwjDkrw3hfeXlY9t79esgFq5Ya3h
yz8DXO7tmwiqg9gC8HxGLLMcxmFpX5Ki9WPymttVWQVCm6DZ4zHAko3iVI+0hd6SgBDdPMznFfgw
OLBy9BryPyS5DWeLEBq0cA+/lxrJB5RtoL2+GmU6I1ZFuaws1tT4Qph+mSFxwUtRiZ7Ly7dHzkUf
9XIN+9Pz17ChAhe9w0ojoXb1NW+ihdapDRgfdVe6vOVFusAO5baQlgk4QZljEGbdSWHFUAE/0xVK
jtsRqzIK/oghPwqoEyfmO5A9+HBrhurIhLawbFOTpP0+aAMVsZtcq22PnfWaWdFyVu2C0psgEsnE
47121DsFPHhzJcntbaa16wwkhHPQJzR2bxmwMUEAHMMJfHYxhHTsN6IkSIVZu69YIJqgxs0/8M5P
PXfmbTx6SKg8hqkC3xFLWkU3O49iNVpif9HWnXVX2UNZb9IbNQDZJ9oecgoJhu+RdlR66B+aQXcK
jQ6xC36W/RADBxGfiobLrb4EjpU6SYd+zpDvL4fgBi4wAUGRMXBOWTGZKoVl+S0nEtNUEjVLzZPm
guaZJSzn2fwstJcP3hZEIN9ZR/DXLPTOqG/H5Uh5mHp1gvaOSz8g/cWo/H717h2XfQLCITR6KltU
C/x+Zwu+Lva8rESUviYo2HLqKHYoJUlzOw6CQZyyOtqInCtzJ1zAzgrINbfjoJheMTucdkPEtwV2
WOWT8mVhWXEKDX3O/6wr9y1dn6wQ7S0RluJBsba0iwKzJcDcj5OyIaEHhs8o0pkt2L33LREVRt3v
Kb9fNYpLsyahEjNCFVyCLUj+Xph5siUxN7PWWj00nBqt/E5Pz9msLRVqkKQI7FFlnKaUPyjpNTGP
QYODNx6T0/MeIehg9dQh+iLZ5z0y9jTNV+dycsrcoTxcg+cV60++DNsxMCAOBPMpjU0L+5aFyOVP
1sCo0rCjc3EYWc2lBwM0g48m+ZToywvNNfa4SuA6F5x7ICEVNDoni4kwZH7UtLUqdO+fj6lwxUOP
gxOPS3PT0n/dzCyYYWY1kwRD4UKxrV+yX3sr2gTcVpGgTn+0swtYNG6bnOkNjqyNujWEE9hBCnyF
WsypRTqhIOcUNhFh3QP0kMID68lVdl442HRVRkdWmtQAttE4N6iH64KQcKDOLxZNpldmC0JYub6v
IkvYLSM+LT38rwg2t/Oi1lboWAQyzo+1QdwZJ27HpGT7/mkrb1GH/mt4Fg+oB6W9gp1ws9WAYA01
qi9j3KPTxC4/3Ad4ehJIMh15w/ZoNyvpZaqp3826UznBpDiYp/rR4e51jpdfK/a1SMJraY7vYNFB
ENyEb2mEmYj+StJzITGWJcTTBNwMYSCMTy4ncPbW2OLlBJW37UZkbqIjCG1+GpFaqMhSlO9Wo1M4
FBXTDkdFjKiKk5Cjh1t1KYcMD+ze9uMzwf+SCiclbq2f6NXpyzb/w8KfhZBwTF1UDkFqe0143Ift
x11oNs6wvuPW/hlO+bdXD9gO3+OmloPMuFp0whj9OgK2VO/i6KYG0WR5DUYeiMW3CZXYFZim+lJJ
P7TN4sUggmf4WjhmkmJdm7hHJZPoBqrAuJlx7i+0//RSO48tOqe9EGJUtBuAaNfVWQudBeo8QN2d
CoFrkuS5srM3ZbzDCww14ofFXjmAUZN0ro1bFN7rpegLP+gkuOV1ByvTa2cxBjZjlJflux9UIajY
z1CNOCYJWRe2O+1q/by4QQxaty6SwIZCRMyckao+qpaHZopteUSxs0Cs3TTENJS3WjHton18KzDb
orzhvv9VkdRJviralhaz7Zks2vHtyLjPQbkEP1kjWM0nrBtC1UrBm5difL4IFxP0uHype0xiSbuT
BOd55YpqvZsYxaNeHDD1i/15IeHplUlGRdixMw31EQXPCiuYBTEGSrRB2wNZOP+xK08K2SLaKNSV
BfQKSNSSYuhmRvCX7G6GV+QrOYt1YeFvAfMorDPShJjOfpudYqqyf3SUw18wwqdl6mFYiOeswQSu
Cz74KoHTGLRxhkKi0c8A/TyvMVNNBOXNB3iSq3DqCBa8eUSTdaOkSY40p1zVJHOrO8QpKwf5zC/H
ipQoWwQCoBwKglGdReOIOfQ4uPk/aQMSesvyqnSyTs42wqhx94SJm8fpUujfmWWMhPRsQjyANMRC
oDnTGjv/X/lpPCLXSVr4SVswbzRjpV65bjWfEPNpW/Vncw6vUgSTTBqNFsn/Jt39CV/G1H9JZeeL
wLX9aKo8vTonhoM8TXnFZn4PWm44eb/tPcSi/FYS/jtOnKXLn1mWp7yn3I3AVecgYDYdmFTTZI32
zobUUw2DXCh2JWow6sZobEY7YgEdB69azSG1UFvn1QW3Kg0RMPWIAIj82HoiLawgzKYf7J78Jeh7
BsGDVszn8Uq4w4Gp9aIAQCDiL22L2Mv8BpG+zlqpDhN6u41KDkLdIn+8OnSqO8VoinbQC9OLXbyi
JD16AHcBJmuV80L4Qvik7uGjCPIMvM8MdiQp/5NfuVcbvAaR2dbhlcxnKIE5c2o11dD8kd1VQUQ0
5zShkIhz2MZ0fFcf/2LWADo934aOA+3Dk8cCL2yas91UosASq/m0ea48oEZXGzj69fZYnXjEOtdx
fGcSdZQH5IeH4F3WkN9B9SCnaLG2FTBzg/VEbINnzxSqzIysPOKyBBfHg5os9+qOqYeamPBg9BK8
S210phhhCdjvjimE6ugtl2w5SdMZkhQDPfVGpJWzfX4YuRRLXvtrXP7P4pympmLhQHLMw6qYDCxJ
o5o8umc71ZxcKZYKm1HQ/KO2R4HULQOYmlvuFJjX4kiDDQZcAP3nb9iii+r72fiAHshDMANmNKVy
I5osSMobTOB84wfoeO8cNMNwFMwOl2HJcarh2duUzN3a8TPULRLb7cglDH0zIyVlJSwxw/7nvBt9
+MFcu16X6AbJwS+q6NIwVHnaao5ys3fbXQLbb4YEbfeCMj7fAPR/mGrgCZMVqsuG5Ff8Y3eBVlYF
2cAUb6RoAnkB8vhYYnMLsxAwV/ebQM9b6JV1cjnDn3zZzKQ7DQhDOgADaSOG2CjHZt35n/kJFfbA
a6mcP1jfa5YqRr+wpbQrSn3mUNzef/4v05rcyHSpxPR/A30m7xKQYnnGyUQAoam49ncLGGBTsTev
Dugw54F10pJ+WWDnZX7f3XW/QPqzijaZrTZoBdg9zwebORWnw92a3KL+8WZPrP5TZmsRM++NtqYG
SO6CkGlnE6jeEfx+A1JaBCyyiSVy5fD8cjQxuTBBr4LGCYG3TfPmS34vPCxNcWYcvXxEZ55kdA9F
AqScpzcO5h6fZA7CjcueyDwGC7yA99n1xv9EfrVS2DPs7a+D0DsC+H5lqDw8C873veMBc/6Jt6ZW
ctdfvxIgj8P0jtx7fevLs9fsls/5a/TTmJODGDi58yo8UKVk5GuaZK/anUXLZ8FYVC3wZEyLY2BX
UXfve37y5kJzUDZIltStI24YY3GfF/rVP60c0bGlPJRRQNLDnbty0eeG4xbHgA5a4JV8Eawecudo
aUwM9aWHaM7hWabpFD9r97PRA1m6ToCPdV8PZu29g+Abjzmwng+3JPwOtffWpQworw6dlOQpgCDc
hkvvLNTdtTQkYbUmXVDvoxhmmPZ3aNrgD0X7kDqaim14Z0XtaFdb8AU1H+UWJoOib+Z/VPDPC7y3
7GqiYOnAMdJRf8ZF2qssSiX5mnvOX93BR+w9wzb4WRj6wY1OpoQUUgeia4cO/r1evTFJ/Hwcg3x1
9SO7fOYn4JKp5lLHr5ByiNcNgfiRjcu1YzHCagyS92Xu5MWaTbMx/nGOlmSHxvwRHRLoyFGIx+ns
tI8BRc8xJB8bBW3jFvb/5dCRVGSX2BHALoGu6tUTUDeSKMoZG2ybUsZ++8PLRUt3ose4wIlmzsh4
sM+MoVtPdbrqYFgjXTV/F+ZFDNGXAU2XWFba5paPMqiHv65ZUtR+zWnojj4miOyADlvVKUgQDKWL
axqxi66EXtRTMc/hRE/WA7uUriqaU/oAJzm9vePeklD1MLGIi2i9FFnTkxFdjTcuzqZkNqes91Zi
Pd4Ir13MSotfpPrFCW1K85KuPbU3jS/SyL06yl2Ci3U05YoaqsR27vSU5XbyjauSUGCRlCYLThDX
vKRjC7nxgIMvPdgzXyN/hGC3dLLEvkeLE66VhaVlwqavyfnSioZAVgwd/ZVQtEzoeQDQK0MqLy4K
aNc7c8GNayAsUXiWhrtMBQGdtVmNgXZq0NXI0U+chE9bNYjzYNMSaTQz2JHWuHiCvj1IDO69sisP
KziySJ71PnlQXgrrXK1xpAM17B6JUMVWnp+Wr+aqWjVgQq1bOyG2nFOMIdwyVcnTq8RBbzJDxwqe
ofyvJmpJgJ2Mg0ooIy34DnebeyNSPSIGW8Fw98sdYv7QXcyObiPBQYZMdcVFT/bwMMdUSuP12mz4
spraz2jMYUsVfI9+Wf/gZod+fE1Kxdk7I19Gbm15+jR/PkWhhb0wvTrs7+vJfuUmNIxHHbujlEuK
BQOk8Qgfn58cASotePy5IEt01GNv14eB/Xkgm/PUT4B43GksRQdN0Ot3cST+t3qZ00wHWs8fZXRx
XWj4Q3xE3Uz1eDOLIshsclPlOhroVHAOZ21NNpAveqMzPo8gHMG9U61RDvt7yG+zW1vC8iOB3RGl
nfIa77GPO6dZlG2cku7atCmkOgITqZRmtZnjzMDZg/GGybufSnWF7wUEvsvFX1SxxWNWLw6qUtGD
ptSYg6u1luGgMfDApowlwbGeQNIe4rRJlDcZAhlSUhAjsydztcL5X1tffbKn3Z3SJsOzLTq7lNIv
SJDpNv+cC3ioxQOh16c2zMITgWRoUN0/vvXRpt/VBuqbpygD0G+fF0oc3A9aCBf+L8e2sS1AakEl
UC/8eI4y2wAWPW3607bwvYl+N8unuOH9Bp7zBfmQBl+IlwsTO62zC97dZUWv47m38RRyzXbOLkyB
5F4DHAfv39E9i+kl9Tp1TkEisn16dHjvqxq+exNDCioNh4wQMBSuHwz5MKK13x0oRnAJuF29swYa
t9zBGvf7IePqFBCSTAVLrrLkBtXFZfy3HrKq13p28Px4eQSu9fPc0Hrz0TJJyT480eeisGAeqEeF
cWf3BY54HB4/da9qM4/VpdeKkPi8hhIh42ywWFIhNzR3TmpAV43JCSsJHpbBBzeGlzUPvdx2hDpX
i22kNbvmXHNets3AyMrCvKqrlqZU+5ZrfhIDZRGIh4I4qO6WueVr12VKigJTn/eLDbPdH4+78Ieg
ux8B3FAwJec7mQWRoz0eWlyc3c9NnHqnuRuykSi15VqwFYNchkG9BalhBugTjTgzl681CWYtaIiY
r5juMHKqHw4dYCfiR+rHQ+GZZC6U6W0iOkjtwZpnzv9oHKQ4xfv5aDtgBVUhTcma0wmms+p9HrmB
3BajzFuHXfpZWbNem+gVAhkHbfrSJ2jaTGGXi6DcLw6qRv4gtwMFLcoGFbDErXMrPdepXQCpJL5v
dQh4T2uaDtKnafPbZlINAPV1lUCq5zGfKWXpARJURIF2ie4okTwtRSRRGppqYD6qVeNMacOAra4c
QrYpjJp2c37c79f6FkrKAyLRcseEH6bxVtMxgWDNuueyUxsZ7ZBqJbOV2B2E/ihacB0H9bCp7FFh
pFnsU0ngcnTsM3IxR7v6HO6PClH8HnsfLSOACSZQ75RZ18cuq43VWFy3PM8eZAbVtiUXres3XWv9
iXRRz7JqdoL0BAgNJ8V/H2DyvQrPq5woh6ekQAD5czLVH/sXsqRvXP0AUMJgtklT227k5EfKLTOn
v3wWM/dAyKqIyDDniLwqz9Sgoblf7Pod78gjxTE7Y5NvbzaxlsTlLbHBLSWWYxSMpOwGqOqFNboT
866g0C6iPN0gXTV0xSBtO60r1w4jcthl1JAwUjQ4rJ2sbSzouwBo8x/0Yd/8VOnK5WM/sDidSX7G
vgvF0XdbHzYapqFmKavyQ02Sa4iygTZT6tVLZM91OAiNJIQwPHyZ13/mVaC99LCsdHo40TC5CXKZ
S5L4TD7g5Y0SSyJjwL2BSUfAXKMzaQc937P7X4n9rEZEZak5/wp44hyJUgSFNPhNI0JPHmfv1ogq
Lfxc/zdjCBgudZ9/98pI8AedcIEoKgn7ZvqUN3blIeeejsSZVokRV9x+u8rtVnQJcBSad2PsKsS4
QJvqIjrQWyXlAhMZKQpi2K/1tJpht+KZkRb56Kk+9PdKx0O4WfBBumjxxgRB5o5V+BKdvxz3zFLB
dN/nmGrvzZyc34b+uX1wtJwCjuXZZ4k4oipf9DojklRYkBgPnsJjheXDodRNtkRAyrTivx2rNCsO
LaXncXlHRT6cUs97+EsVPTeIk1I7lBpwJvomiZQkE3JumYaAX3ziTcGoJ6/LZN7ECQqAZLUFGp/p
NY4/R8Q4dK9OZZWspUTMAgNRPqJQGkEB6imqka2qzbYmIk965dy3RcoUte12287doOBXoobdqWye
fE7+ZXHV/eAqRWjU2HteSwEWcX5g3Yu6/S2jsTi0qI4f4NkCxAv3FA/m7cBEkkQFIVsbxZ3MZ3MG
zm5lUcqNrfJFuV2EcFdZRDArkwyeZY/T+dg6u+JEXykSZznjeomARXVsZpviKmWVhgFAR1vJ1Nt2
MwNOdx9zwKGFsVoWoEd1ezESQm7vaTFq1msppfXCr+WiMS/Hq7Ummz420YZmfCxcnfFIwOF6RkmT
Sl6lL1xlPUUhlZNFwK1xUabSGjNz11HvSMT+6SxOBnlshKq6dLwMWl0x7EWnZr5o/YUaC6MRdnfc
PdnPy+pU1pVChWqWdfp3CcDQYOM//xPQ4R4JWMBW7G67kjhiDG819RgcNzk0/LVpoV9DZ2yI4xH3
gQm5Hk42zhx1oWCEKgh+KYCEOcO7mDEZFaOc2wXmcghe3B1HdJvkJRs8ng6MI68JwReGM/BIdO1J
wHFjUYBTOPWcVdnoNTR+pVc7B8CuBzqz8Rrl5Yn4cvjSw8D8ykQHWjGcMWyNTl6gKwrWBqJloCyb
YuJAooFGxnz7CAyf07SBORCt3lI5TkjUdA7NPHNNQ4M9tzX1WXO+YDIlsulnuyPDzwHWyCTlTV2j
jp1iYkt1P08iyop3R/jxMvaFcvl6H2XnTr3jWEwZkFDzfhyYGBB1wyHOPUIi2GcLPA0J2RrBxWoE
/5KD/k5fcLFGrQO5jz92AFKHaPbODVKBNLyzPM6FGdbvsgII+E9afZmpGOitu8SZQ813+8ApKQ+n
CISW3h058mGF4hy+PDJwO5jxux1t1Ca3zmDOlOBJ+zE1EjFIQGyJbHzFeS58ZI7JWmIGCr1FRezC
im20lHkl/mEqUBn6vHuAvRIEKMmnbh7L7gz9e5jZige5ZxKzOO6Wcu6NFB3q60zbeHrQ8vWISwWu
kBZ0fa17wxlU3aZ+WvosLPRSeQhF1yDToQqOAhrRA2rKJZPKLPGpx28X7Z1RgHm/COJwiIsGlasA
tK29E7QICDtXub63yVtGbO0C0CNgNk72iLTzbQuHUowuE7tvkRJ4ibyG9NspeRjGLB59EW/QkhCY
OkKi5CB87ywNMXL6L6x1fbqDmOHreKp9j4vxGGk98D43KJ7s7z0s0ad1uyLcRwvcUYT3MclaPmzj
9DMcLHu4pMLpApdHJPD8Y7nlO8N5miAREnJh2p+F98z/AzqS03LXpTemfex2X/rPRgC++k3/1f+E
7VUAqtGIE+HZ4HMzEpfJOta0mrmxSkNMMZ6B1kw0DGlEw3qt0Jqly5eqzY7Nm/NkBue/zTKvgs+r
4RHMujAbxuf2ciwqO6wb/MwNSr6I8Ra03pzR7q635sLVKbpdgYjNVLlUZQaFIozUkGLIx5/gRPdv
2g5BjIjZblYze8Q7azTIOerz5TGwdb6BUViEsqWozmM7saTAL3aSFIRTQ35ljkLoPeL4QK8T00Jt
dFHXe78RKadg/TtsKBGEXbI7Ns8PpYZ8nDLAhWTnOnJWsckWHoGyB4gELDfpNkTPANr9BNRkAyiN
fiuUYVKL2eFHvfuKVSF3GA7AbMRZ0/zp08VPQ1R+14XSHRcyYvZr+IJQcKyNTHBTXS22iKl4JDSO
0esKSXZ1XZdpG6/1ImCZxkPiqAOsudHL/Nf8Gb8T+bmUbEdjwb/jptDKVjWVR6WkEn2D/eSsISqf
EZF9/1O9seENWP9LiZYxInCKJSg2J0uOrNNtD6QRnxrqpU7ojvMtNjxJITxavrDTan2MBD8dfYbQ
ILTVwIVhqaCYJ9GT9uGCXWDRfNEoMgvtWiE63ySwu1PMH+yPmUyPr1rVRWZUyCsJmh8nRSO5GZoS
eqZPoan8HosYijjnflcmYzvAYDXD+Hkp13wk+C9th7Is7cwh1Hw5cFy/leufaKOTrlHhGp6Tivgk
KTqZMa4SPoWGK0C0w8MpVZKett1lpDhVbrmJkPLAixIYgeAjyi0SE4pXZpBmXj1CPzcG7bJzbPKH
rHC1cD+MMYTQ5NKXRSMTg26wS5vPeetAW1hReKt8beJMBtwHZoJD0/gweYdGLByIQQ/I13rB7TOz
8Un1RVZDPJvVI+JH8B+0RrZ/Eb0HC6r8sa771EjsfMFHfBm+gMlXiJrni41v+LrXg39NNvwrV2N4
4HsiwNVs+QpF1+L0JvyuaodcfalWVPVQdCiRqDWaoNwnLSSB2b4vT13ryFbLpFR9FUx4Rz6kdh63
0zsJWT0YNHgFQXuIl2jLPn7hJDPk8qHgBP9pWY3ivBWrTCfBylyLP+xJ6IpylCxec8oaToDwmZ5s
EOVtC4kiUQ7EFMtKn0dbfjJGuchDTwr0KQUnKxXNPLNsxPx0C/55jtmnwF319dyNjQ81BV4/jezX
f1OfEoT1jbDJMuQOZqs2ffFfFXozXTcsCUaonMNo/efsPVdv2QI/HeUDmg4U/5zZWocKiL1Hwv1p
NPinIVhh0Cn0CWeseGlASLLZTh5Iwrutwhsch1XwAH3k5HVhFzs74HbGoUsTZBS8BLtRpNQJbs0J
Kk8pR1W08Cztxu8X9cJ+aFQZdV5QVDKZVBesN8ngFcNemzd7RcCGJFn5CGKGZbHIn1rRQIjSmiQp
CT4TQKK6ywCaQpJwTA3DwTnBx0qd2p6teegaBphyLa+3N8weOHFskvGBX8CJTtDpAylIEs/jinlC
RwxXt2kuR7aDcVYKnCJHigNYSrTN03LdiUtbACe8oDbTCmQZG40bWD/NPTocr81cGbm0Q2WUbzqT
akJRBtq31eBFfKJ7s9qOg0J1oh+fXLyXhGAXRP4PURGFUfUAXCBJW7kwzPWWx1u4JMItKXA3wDPB
D1HhxsLug8hH/MFnQNA2iOdwKvsN7WN3PxNaQmKO48ZXmuht5FIv2F2CcH2/W2t2Pflbud7WZyuf
HUdmuU6s04rnFSTlr6NtQHdXlwbiadJdPpavl5uo5y8cVHzKK1335prInBnEa9JezHoWwM96S4dY
RCzCHI29nQwyeLYM0HmP/Cqrya+v0zbWTm0euBGD6UB5wrcfYdy+TWNvaHq2DbzQ2zRnY8fHopJV
4nspZgcrlgaPs1H6o21NWKVmamu+M/nGudNkFUHHcuHJKYvZP03YAMBhg6d9UvMGXE4qtQmnFaR1
gJNFG35Hhy5z2Jv7GinTibj9lW95Iww+HI+KBKjJdAtzR8SJCRyn6An4MUrBBR0yGp8eosUSj3zl
NRdCRN6QT4GkMR5p47iNfJNLdKFa+oq/4Iw3PsjKOIfVtXNZMi8Qi6tYuhd4ZPqBOF9BbEB6r7Oc
RcXL8yhzFGRUWG+F6hdfl7feRGy8pij1XsHYs+FvgXs2nSZSEEEwLIEZNEBm/dl6Abw+zuAb2cXU
JkyvDkz7h4gt0UOHdAvlpdF2NChHNMQSQS47scnMEkryDgkPRUtenjC5tOPGQc81C/5lZsG09axX
QQgAMk1WvPxk56sKejiWJ4bt0hYW2ngqbcsZ0sFWRHxhKWOXhqoTuU+dfD8r4NdAjBUaVNWT8lBc
ea5BTado+aiHwR1TWDHbN7oU3eCcHFu75g8xwbKO5W7k120xV/hWJGiYikrdFDh6pb8P9Ya5MhQI
+xGi7ANxqg1iYuDExwZDkD3CjQa7pslS0onSotRnhKcBmPgBrcDs0hthoq8OOtv36+6/hUrI/vXY
SuvoZ3Jw7YeXnf63a207BLa4MxDP9UXcUL5rgoIKBSJQnq+ScRyQWx3P74f6zsS8qor6B+z+tlW/
+4RiFjo5j4By71l1kh6BAxY4U4tnRwu/xrFXhHgk/BtvktgRoFICg9j9r4XbidMttPz9t+xkgLhn
btaOegyGocbX4BdJlPYB83iBthej1fRjYOfCz/NPNR+kN/MjaCiqjlC5+R6xXT/9QwMCdyzGpulX
f9Lr233i+JtEnIhcQeznXK1MixNJbPPruXcPUedJGvD45GwXG0N36uDMSSOjr+XdeJRn6Tusnrkc
j/KJwLOC4e/d/kLrEUyuf9ZKseLPVyxuMWry0Qdh2yf+Uotdwzx8hD+Hh//ZZO4xSsnArOqcXdLF
IDA5Opqz4pQ5Cr2i1l9jY6W8NjTMcKWu6XYQy0NJVTqOOPo29ezQteB+I0JgooojClg9NRZNF0Vr
q3qKrCpwiXkSWJH6z562dEQh/N1+oX2ZDRHi7oNsqqoruFhS02c/1GStfx3/QGh9cxKlr9GpjTdz
XfH77JrnL/t0112I/dvc/iANGSRxtdxEJ/SfAhhXlNgDlu+sSO14F47vpXfubomm6WYpStPzY76v
63Q1RDtJ41SV2cJc9Qq5LKHh5OXCFmntBzx/OpTmNjwY0vzEmFGNfbAtx3cJm3uvWjK5UmkhTAeQ
ZRV3FjouF3fl8gxNRIZhvdfKtrDZRl0zilRs1ER8Yo6yidYDuh5fVhlYEyiQ2QT2yS8+SZjbHlmd
Rvs7WBbBDB8U27fOVEkCpOv+V+sZ1o1yTQ0ESxujqGBbH+9y6QCmXeNB8RpuVndpUUXXrWRO+0EU
zUXjkjIYq0ANuruRWVmqNQlNhw9aKVLK76aNKcin0gMMbhWXHbiWnbL1YJDDs50fvFHLTg3LAOLX
Nt3gBbUxO02Ditm2PWIkLM4AJPdgFxKB2MW9BxQY6hrhdO56n3+skbIGoq0jU75DfiLWpgvwgZpf
75xroBpmtb5gLGXC0aHUmAGZjpt82XkGFhk/yZjojCbWTHiZFez/qeW5sfNv4cd7akyJQs6PcpC1
OjM+wxAN6Emg3oRgXOMl7lI/UMdJ4nzDBxPz/oUQ7aC++kGVDEv/ffzaFNdvwZISbfJAxWj3u5FO
hWTXNnDqPSljN5VyJFvAu35i4NzJpWFF63I8y8+kOrsmgUaJOta+GvNvYYoGp1CDHeTQiOSB2cI6
2GddH7c93b2epew2yASQg3AVSin0vEo+CB2X4EdP/NG0nHNqIL/HHSZTJHrRUMCCJtbbs9ISnVXO
bmNDgIBU4/ZqFkHvuC6SE4+sUIBHYn9J6Ce0o4/U25tfjRzapjRk/T5GpJXZ+qN7e0bWDV4DcwXS
MH3BYlwnsqh57DUdIf1tPqbHCbnBFjT8VMP3iOarAO7DzpwjoTeZuAK/KWrjxgnWcLAF48OylZIx
Ir7LcR8i7hHZ1LElAfDVDS6KmFGKqEC7extjclwJ/pn0NLXps8O1uHFlO+pUDAxGmTQXebB2hNyL
SJEcIe/H0U8uhyyaAn+XRt03sSI4zKj+xrDEUn8BrCs63pC8jjVpGQEiwVvYe41L+dCeX3u2zEsm
3HXDumKCCp2ycEHLZLba9Oi1OgcWVRS9El4qr9g1W22+jsg0AkL5Ecl7g6syixxSfPABjgj0TndQ
xOYg/3Y12HQR3HgDFA7ZpjhxX5HTymR3dX7wpazFQwdwXxAO5p8R9lVwKiMj2/L2xqBwYmlPo9eR
zU20nyfza7gi6gUqUHu8+EniXgoa9d2Xu0WGUBy+rsQER0FSkVosNJbzkTUjOQXP9Ons6tBQ3HAW
mBSQSxVja9euIF46dC03gCXREZkDRFXTLgagElEZ6sfSmt0hkUNUSjodRzr9niZwmsrTK22YTpse
fh5v/1HPnPthgIZPai4TyhHI3lysC8hfntAfLv1OjC9sGmuZ1oxaxLSWXXQLstV1oV0D+VrwrYGS
CkErdlMlA9uSF1xfa7ILMhz3GpHdFaZDB7hI9z0d31F+MzDzr9mxV0X5vWvpfByn6beSMh+DUsnJ
Kyr8cl9mgh5U31AufulV/hRt5JgVuv3iZ5SG2lylYwHt5g0KxMBS7grUqT85yhwOhLH7UHucxX9c
iCd/XlYio0heYGJzankBc2UUt4MWtERvkvVWnmT9Ukw+oH5yU9vhhCor8e68wJHKfIIcGasa8Rnn
rueqVo2MZg55XCIDhOox51mWDPOFxexLJ5Gc06LrcpOzNyeoK8I779lTykKSGe5S8JeB4DWnCq/D
1KFuKYq7gKW8TjqbhEW5e+8FoXqWlBNOO8do3WRuZUvl1Tavx3DRCgmcfg4q+DmlBb0JxRT9GC3+
90Dpjn7mhDh+UiUeS3wCT3kjBXGAonuC9111YYRf1fH/CEbMS1LDEum3pSSs2Ou2iH4GShwUG1yK
FU/EcG6eqC403Iv6UNVbTQUToGury/AtfzCZfy7BMHOyH6xiWpnpmXkkhSz0eVVkdQaDlNvXRPIY
f0nsmfrFJZZ4PW+pDBwUqQxq3ISFSjcBnpgmw4uluS4cfviADf4Wf+WsjkTnZaUdO5Aian91wPe7
OWX/qzRGJiL2OF7CRV3+jZzamtdpwoZZWtty+/Whf3IJQN/V4zd8FRN8SrJC2fAF7VEuOLoF8Chn
ankXsDJsJ+QSyDs2t64iaf8K1v2nFmZSf27p/NPCS9h+u51wbdn6ItOYGlVMFE//Ur5Tr8m8sRzC
zxovsD+DrdJAflclIA30sAa8zd4Ju1+/7v8dFUEq8AKDG4mUnMUDJ9mJsbIowmRBbtj9MXqZwuYJ
eHJGZ5x0SZUanZLuMVhN3qb0mB+3FqtG/xahRFqWlbh9QgJh9VQPur0P/Mca6Lu6JhbKHI8BSnLO
yIDYvm5LleIwhAZrQ1m6CO/SNx/bFngWGKxN4IB8ZItJw4PWny+j9mDiYkhJ7xUj/GN1b2DoQJE4
16G7cDuj3qfp4/jPcnvlyKuj21fReA9dGJgzcvS8r1JAOxCpV/gQH7PefyqLluBIWfjnzoYvgQeQ
SDn/pSta0SDWkMVTR7zdb4YDsaGQjEX2LGlVZgRgbWeTz9qXx4t4u8w2TcEQwkty366t9Vl4F3Fr
1YXHy1sl7m7cV9nv02yOeiDZyz64NdRWo6PgiGi4jjIoXLCBsD42uqQk2AqWw+1Gcy4VywWl9FNu
+vdUCzg3BUxMmpZocWTg7gKq0zr2eFKf8RZ2FTYY0NxmTSNkk4KWmev/e1YcRFxc9iysIrkL+2kb
5CtTNenjQKZZs5ozEniALdi+CU9wfbMcR5Q75lIurNNIuJmolVsvEafDGxeBWUlvwOiSKYBqbB9t
trAeWZ0TK+4c+6QB+TwxSmQX7BPpLa5dPlbMP+iJUZ5Iv3zEB32qAhQg3NA/Y501Wj2rEW6iDSRy
WCuIAC4Bre3c3IMpX5+NYeNd3RVBGeDu+xTj90vFpGzU5GhFy6mcsYDnubSNW5o7cdquAv7i1noJ
fTeqMT4zHr9O3l46GUGPgEQBP8o2OC0hsShySwNYs26dBlIA0d4gZ2aokCE61ut0h35oYdZf414k
xE6sNACAz+SaszDvsOoSSTSQzFUlAvcQGmEN/MT4+l5gvuJOFmI/CM+WKJLxT3rXCwnbzaDaNxnd
6h/NJ2QISDc3xAQ/3JoB9S+kFHEZ9gFMYjR+Z8LXdb4a/5JT8BSYlSyLBvjbvMxH6U1zE6Jz7QgP
c+1embRNh/raDR7NYbFEjldb91b8TlhiZ+kUmDEZZF1cokl+p8VWihF2wN1A51EyZPlrmIHvEipR
1dIYr0UB/ytI5Bkeo8u1Rf9EiXWodwXiHkUp6ttdtigmbdzcek1UXmwXUFQD6DJveoXtG24QYDo/
A01/R0/d96CXdcCe4lVaSVZZ35uX5hRRdbUxXJDOA0O9P63E5X1G5MY/TnQaEXG14iSMWFUh1FM6
meU3v36+J/Sgoi820PD0lIlgvvHUVbhrEvA0PLG1mvmy3xxUoVEkxprNbuR1bIlTn4ZaQYqstI2D
a3IE/Kwco8J4uNcZlhCnla0vT3sPyoZ1rDT+KIXQJjFRGdkyLZY8ELmu2o6eii91ATnQZPPrGyMg
l1+ZmV8qlp63q/NarOsWndkkwadyFg/Lh14cPuMTP60D46Xnram03ctid+t9Ui14B5t+/Xu/0HK3
6IUMldoatkLJQ4rBMOrF/U4loKVdPHhU/sl8AFOiiIRnfzAFClMElkftP3KFR+bzW15Ef0fA7jua
t21cDJTO2YHZfVeVK+yIc4hsV1JcYCL47cGfrckM1+uCBlcqn8pt5N7/KrBEyTO6j2G+xM4tYFpa
yjTX5WmKnzGNTa/4jzpHem7TDaRAukOIhwbgAxm05+elpmkykaBpKW5CyRd0RpRkKVlWr9uiJQJ7
BlSowRUSXZ93gGz9RDvx0CThIIxirEfIbHhA4dEmJfNFZoq1WWyG2I61LWRYDGLVPc6guTH9+GSJ
hkDajCSA1hhicn8JbDQ5k9ujHA6PetD0U3oXL1JhfWTgF33+JVE5INWPrzEZ/7Z/D88Noh9HgLOV
0BOe9He1YDFlkd2OXN3UKCjLYI9lF1XW6pg3QSb1cH2SdUj1RySkQAeYWuqSJ8wYDmP1qm/oz0jk
y7ng6KSuoyJlsw2LByQ80IZSavbjp5aTTNvnX/8OuQuErVRmB0SEu1VnohWPuahVnYF3+EWoJzoG
sknRMmg2Z19404wJxenE54Rbw/TMK9Qk/q1Xzg1jOj+Bs6bPnf6uQks5uJIRBP4kGIlEwwYxEF/i
UfUgqu+MjgJt3DsWATwdJGgFJpRgYjcKDtTi0rf1YiDdOdFR5GKcAbFpR7VTMMT+vfyAtY+CjgsJ
IaFs33d+5NIDQPKsqZ7q9CFJN4ZUVpgk9I8GBgjXaRDlboI/kloAIrp4dVB5heAYQ5CKVaQrwqzM
nS/O62v6pctYtpnxELMF/V+SfKym4SYzW3OpTYsGs23yO6FG2Btfx6kg8YBultFRa7wfy9DU8sa9
ul7ZQ5b1BRiQ8oqRIGQ51la+sV2SIfyf2kTVgKKmpOGdFdZtAdOO0VHYfy+QXVEtWkg7OaUlzZx3
H9SnaOMfVJOZEzeTi4D5WdMj3JfkOzCoG841tOUikQcXqaJ7NoSMSCtOU71GLJ0U0IYQbf/TcGzD
gvfmW1QF/aksyaGKZkSjGg5jCV7NNAWXROuSN4gMwnkAdPKHnG2AcuRXAn+t+ugnjEe+ng5ePWEX
aUZa70hE4ESVM3kL36vUOzBsspMxT789yDa2uY0u6J1LLFWSfI6T3zYa1kf39DMqD0b3xhNHNTiQ
HzokZwxewKHkXyL3M2N25MhNz9goH18fkpoZgetshs7HIEnxWiIs/PDIMAkkgr5jqwPW6qZZS6Ey
RSNlRvc4zeXUNce2EXiSFbQl3OU8eLP+9BqZiAObod2856bpS2loAnulDev4dOQR6BxE9kY86ElZ
3Fl/iaYKndRv6hnHX8nu1oYDiaV3ia+82ZewBzqD6BW6GcU8tU20code3zIeXRDDuvGS0aGLIB9f
YwzXt/EqOnglvUPpcXy71u+Dm6iqz8Gu8bhb9wAigmOSgd7LSkBJpaDizLenxwlrcDzp6PGfKntX
g81o7/bs4UkOUfVFLbwZ/jcJtfSYXVIqiCRZDINq2PKVCaPMqw1+yRO9WC47AYBf6HIfCZyRWE9n
9+2n1kmZzZOXW0j8xXBWMiF1Mapf63inBJqG7Saz81+LgPw918QChGvIv/x73ikWtPiazi6hA4d7
knORpPu1bwxsQaqAIN5PqvdoJqMzzetRn9k3lGlRX4Ej9QwyG+K7Mwyz7C5NVByyXywt120u/ViD
WIox8E24gcaB/FueqgYB2PWmjUpn07wubnjmnZ1TgScFSDobuJtH2ViorZ0TbIkLOqH5YjBbsE0x
1cLDNjhwi7np2bOj9rMhphkE+exioEW4pJ/2UOeYGJBj+SI8sIxr0yz+L1GD1SvoPqMy80mTBkWQ
p0zXkGSaIr6PCVvvvfrGYtI15aetx+czAHcYHrXxUVEafXVZN/QtEmc0qBnhYnOgw+6sWkFESlKI
gs8BqurAvJl3X1lX3WzAg5IdC0/QLrZbXQKhwubHEasE2zstT+Tbq5/nTYtPssB/9OsNNes/ZXgY
3NoAdYFTAsocdCXJ5VrNn47KX1h6m0plha9vMGiy7YzujnKpoZW2NZu1uRmrTEt5Rl1SnXqa0tJ1
nnftsuaPsnWTeNzs75PrqHGFFbfm0ac4J+DcVsXqskozt76KdKDaVO4GzNFvQfXKhNQsLO0P3DBz
/V5hj9T2/SyDrHAaH29S25yjMxl/nDZUJFe+JQL2/2DPZjmOA4XnQYwmAYS1FYMkrrmJcmU0lna4
3wSwOollC3sPyIW6QJeI4iY1wQ0EgbhwxWqRAmLYVV2LzikynI9IsZnO+GrfqbhgktUHRqstxfRb
2AJhTV04LReI66pqsPXA0po+wWg+24mgyv/7E9Ut915p08swXzNfYi3PEj+fZ3gAzCyzi51JUR87
sIfMuswdFZvDl4qPkt+lD05HLRhlwHuptvDq2NCTDHatKlsOxnymvbPUhjqV57pUiQU6dbc0g1qE
HzL9NfAb1luf62unkzXMe/dZNlm6P2SQ7VHBW+/AKK3Hz+PJ8dXKuK6SM2vbHXdfv/GZJfgMys1a
gGpLuHdfX59Gwtc3ctNT/8jZyY3FOIIgZZMwAeE12tJBeCDAc8v3q3XYJp8WLro1XneTu+kfjs22
i1XUzvLyyK6hb+LYZQTtQza/TfpME2a6HhAVOXcMLUfvyPTaRE1l0j/csbiIIy8ACrUIsvM/sxZV
ubt6IzmD2cfrT49SyiYQZRUYDdhRVIVoNjvVTmryvGcHrGEZbGz7W/muN5N6yb0jE1NVNEmfXNdG
xXl5FBUlF5UtWdepRu9b8PvUkF2bPDDZ9CH1qeb/SZl2UrM3W5DjYqvCn5WfVR9CzXA4ZXXb1u6o
9sT8AdAx3Owb0qo92D7gqaeseFCSl6tNrJ3O2ZJ2oTf1ulWFpJly+L/vOep2hPgaEy3Ct0B9//Bl
8BOQekvh+Hvqpi5u2ilo9shJ2RVJhiHuVKEq/TP+IoeU+ctc8n++krhivrLymlTxCGAUWe8ixSgO
qR6GfXnmuhsRqDrofbiA83+LmS5RjFzQ/q+EAgFseCrMeO8pzFRFkffZvb3dfOn06zWRqFKKgXdx
VZLIHkeSZsHYODGddaKYuvMzNEiV1I0G6PPMfrNyMmCzZEyX7KKpqNqPftIS9j2lIRQfywbNrUu6
FiVfiZ31/C3wZRppgYTYlgcp3DPy1OgopiRn3quRC/pcLpEaIVEu+iwUdAmbI4TFQMH59kS0G1+g
XqU/a7Fy1Lde5r09gqfilMtiH4SjH9FluDZ2oo7nEPFBeCGZXHFzlH5nT7FCj9rcL2PAPbzm+gFz
xWmwMuvmVKTdfu/lL5/XwGmVtVzcQwu0u1f79lEkyw91LPNaG58w9/BO3/GketV5q73uFTQRukd6
rEDY44z2cR/VL0OtEXIWjt9rRNIhE9ViVvEXRPnlyRHiw0PfqBHF2JR73Q8vwGn7eVxrgOBUfqnq
DhfHIrNmqc/yfyGY0ib70NPx8awzJ+UaaPkB2WNqONEVe/Sa8YQ7iUeXc/939lMIwbnzeaEIUHji
0QnAiRWaiqA9Wn7al9o9tZt//wMOvCXqb+lGiBzNEoKcJCRh8k/4mp9PIWKv48d+jVAHqg4q0txH
4Ev69J8MWYBrj5izRGrFVB/YZK7wh9U/1tsVkaL3BhXOfRZCFk/MixhkCk+paRATE6gPgoaz+yvV
a5H6Hf0D9ukuNI9Z4h8E1jYu7a9leOePA0Rq+d0SNV0QDoJBN2ZcVQCHvb9WHOkoT6eWWabj2+SL
oCyeaFR61UrzOS2SKKYoftgNlDTGPAqCGYgEOBJDQmWx8HEpAk8rC+253jOfQbLGH/FIGchqbO64
pDaXgjZ+MTSs/vZUcCVrCoei8Cwt0ZDbGpMWZqEcniakf8H71r5fNda1HfqpzTG6iNnLYegJYLzc
E2CykBdjj9BOcr4kevPPjQkCNj3x9078EMERODqTi0WkW9I4kpYU1NCXHyIBN9WpMislpZNDWDtG
6PirAPaAkjTY9eQ5Y23EnU0/GfHHgY6J8ErAA7giF11PRQU1yuQatuE822ZQJxWal/AL+vFQ90j2
aRU7on1LLSDIpZEDo4q9d6m/4F7cQmvPIYDtlltEFLiIA12nmyp8t3lwXFmECrwNq9W6E/N/XVO3
sXz2zdtvbBJQ+HXaRBRphxnmMVv2TtXp/n6j73nwTO8ZI4AJfg0kZ1Vq63K8IVAdbpso0tUvujEq
VDbnWoDW2xx9qpa79anE6ddizHFokCSFm7sgEPpocBly0MqBh16fC3ZUTTqze8k2CFtCSsUNKiSV
oAD9aAoB57Oih2rtsHhcRkBufURpcnZI51Dka0o+0sov8Prmgrz3r1TYBTSEWY2B8nHceW7FDSHF
W3LYqpHxDH0gJ93VH3+KsdXLWD36Lkgy4amMYhGoaPgnHlK9o6apP0Mc9DiR2qAViMKL2VnE9BTw
ukMJRs9ZZWUFvsLKwa6UVu3SRUoAGwREqWV1n5hGYNPVG+XyjoR38st5g3lxmqUHggEvoj8g5UtY
KyDLV6yb3TQ/z3TzL/10ORX4ZgmUnlEcoO+9r+aQP6R1/TIvlzSADvQ91143HJDF1WFC9XGOPHqT
mUKj7Hco5j1JJChnfxmMfZRS9+wRJ21VcxAMNxoiusdS2h4gqCse9WPgxAJS/InuEHSwCJ/hPlFf
zaTdBP9si3lncHV1F7MYDiejfBtssGA8cwi2yAEm+2kFVMQOhpFLsZGiZL01mYlBOFOsvaRJlAPs
PpmY4quTKew73iO/RjGnYPEGVuk4OvZwLQo5DsdSk6TVFTGC8/Shp+pUgFRFBHWUTRkj60wDlay3
G5g/znsJELz833hhzlvNyuMI+yT7W970mEU6xtn3I0/1XKJ32ghi81vDqZYn43q/5fXvQdai5hDk
/uQPfOQmnZflU7a5/02KXyHYLYH9+XQPDaa0yr+sSaG+HY3IbSwjcEhzOWqkP5Ij5QiGKo0mqUKf
xA806UvAKssWyY6n+ZY+LLJHJ/Vd+cEuWUyTEJKA6Xcd8Nz6SCqDdiZW4cKW1KFzTXXZBnfkdOVq
U2Zk0gEleh/T/rfJxQyHb+JbznbLidombzVyPGAq6qMUI/saTfTSMqLag8exd+8wUg9ODZ3+BB4M
CcUMk93eK5x4WzcZ+FvkzvR+lxo2Yvsdo3w3QPkorxaBNoCF1Ubl6lUi6Da6vRQLoSV5g6J0jqqf
X1aoNN/r3XwcW2a51JsZ7UDytz+OERyt1+zr6JxbQq4mmYRyuowubtWx8MSmBF3I96siSXsXuJDG
MpJGCkD5PNwcdfeGPpdsNkxM1nnuK07l2e6t1W72wATmaSLwZMjfxT1Lfe3VnH4PqF8M1rf8RGvK
xD40ZwMVXgavZ5NcEetpt/8MGy/rJdzy0yO5l+qs84H6DGcIuBXqSmBsTSmytUaT3zdDHKVv4Qba
1yS6/NsWlLlb64OeFjbqdlsdc+Ydm+ZoX86PspRZLO92aNfyyTkUfm8AshMpuSke2CyqhOv29UJk
6WK6Pm0IBOTA3dSNS+DfR5TO6cHaGmt+3MrjFgSHue5hlKjMcyccrXaqxBoTiVwDDhEZTY26Ntwv
JbINoYHaA6Fz0ES95Zx9yhwUpSNwVnONfb4lr/zRBuJn4D/z8MD0ST60GLyZv+7zVZtHJPYGhudk
Axr5ru5kyackCT0sw2ObZ9z/FFv+qnMzpH1B+mqOj2/d67iRXqGK6azt0oezLJYlagrqvsiKT8vk
5VADChAHbHREJTJpULk4qvDLwEEDJk0xW+AQhV5wtxSQLDcCJjWB9766dWIifg2XwcBoIKg1AYoG
m7+4RfC1kU1+7/349NUbAE1l2Qn9hnriJgOgkwey7Lr5UDw2cHSIei3+nQuOq+LUXl8FALWGzmwy
THndg5yjN+W68agidwDEvg50FwrV6jCmD4PNlNRneVAfU4X/R8/32ONIKvjS7fIFOZaxZ24ntbnB
wjQ01MLv0M1Rn3MzjakddBRwmAoySfEBMYwTTDwylPW2qzpOKubmiQ7LZhKTVkPd7cymCEMXnI0M
GXhP6oYiCD6D928eQnXY8s//qFbiUZCSNQ/HD7XlzWze/0SPJHjq6RuJgm7/JxpzaEYkcAM7RQMF
pyy9F4PyHX9DauXYWURWZU/z072m/6JLLaOl0fmwnODW95Vvpb6V90W06B+471QGnnDTkLRg1F6b
o/rYVNu//Q5C2nXfxCgt8eA03WzRklLGPGT0uoSlqoeqiH8ms5x1nq4e+TqO/GxVAGv96TYt4lWL
DFDvVDNNavzTWig94s+un1B9lpdm/rzOyBes3E8McHPkJBrBIDtjadVsIMyg43569jhpKAydTDBH
VUfTMVjgqGH6dX6uMngiTCFsubSiyi7WdEJL21dcVu1/sQY4WgbMElw3GPcXtik9VLSslwGId/5m
6/XEOINNTyQ0oYsKpXURF5J/seJR9s99V/i04BuBzluOFd9M9rNFDXz1yq0MsM9zY8kaHw5lk2IU
oZy/AszTtvU9mKp7olLq5OT4nqyDaNHwOTcbKqaZ7lMe+kEQiUNaoilk3SSSeQQP2n5y77YxfXL3
ZzjM81WLN6qGfOQDxrIeM1qwpxyxER3OmziB4aE1yN7sUzoX1nv2NM5tgi+KOP94iEGCoC5aggeo
rfE2i8D43VVd/vqoC/CLKdkhi6eKFgwSgDPIKM0hcUuYWrircoIO0NFEDZlw1aTMDiRlodu/cslJ
mc6FBS9eKmhtPmWAS2mIuiNJ1fmT/wfRqvMr5lDptYPnFOXVMx+ZC3xQgGncytUf2J65Xddm34sR
rq3OzjYSoFkm4GNX650fTYw9AmzZBPNxOPGmD6AODyux6IJissijxn5oOsxktIu0nrGPyo/+xuHb
/teXT1zTddp9gU6pbE6idpRmh8EUDxdLhin+JF4srQTzP1q/SlmrwHL8WjxTbiT9Nq27G1enA26p
Lu9ynzJgo5pjmMqVEzZ64X/EI5cR/Tbqze8E3qPc/0Fz9PIol73dls8y9UCqnFZYYg+kDBC5Fsjn
N7fKAK6+jDnmetsxE7sR61J1Ms/V09h7bnro/UN8psx95a3ZBv34CzW8nKOMQeCjgdmGinYprlmU
3gA8tkCBPUeEVCFG2njeLGGkn+OeDespY3TLxtnE7DXBUHy8rwM9QCApDTnBgGxefN7V90SRloSA
zCoMTIAFRwq5ZEXvTlVsd+O5grTCMuKtNI+zXCWwZecnOb26ADbu9AaxIujZJTakGYSbyLB9rj2g
XOG5SmnGiIKJWcOWf1zpHADQjmG9bN/bKeIvIuZ7bccLkBik7IeCJQv3WxAdSggLGGHp+X0MoF9J
iYdKiscn9NfUCE7xzKLsdqA17KKPJqNBORFMcF23SKsIxVvPiTcqPRExZiI8HFfykL00Twgctg+f
wyuA/cl04A4n90Sh+IMApfi9a1TIrfvP1C0Wqg0+Jue1d7gEn7xoU4yA8RZ8rcrMpCiv+cx7Tlrf
dJjUQlstG+e13IukqtcADJKpLR2IIQM4MLLoSOg/gmFdVgi97Ar4ZDGwGq+rvw1S71kyIArvUoMy
p/Yw3/ifoT9f8F3LjCGVUYjXtG1zMEDoZcY8X7zuo+4Mai4e1LfFRzkPlCmYPdB+vSzKew10G760
uqW9pUs/W6pMjSAeweBfvi2GSiO3mkRb3Sx+EUuRQk25ceD5uMZIkvO25DVKybP2nTIXsVqSdvPo
6jMHTgJX8hWrbMWB6kW/2eu2r27jx51Y4l1qFGwLlKg9EVJCJIUS+6asUPS5LC+XoS7jjdVgqm22
jXqL+h4tiBU0cj9MUQbg+7eGw9vcc2+dquwhkmoot2ubFDmXcKJKeSp+4oc7vLuN+6sxUrC2pJ2f
xB0ktpmO+3JZNIJ9WqL0Uq+Xu4y/BaVcpBzUQ+EoLIEzHPbTx13Urkfc9L9nGuB8NFraDYvMDHLJ
CvzKj+LyvldHDkpd4jT/jo2+4sRlwBH4JfaQgpyMFGx5i5PS7dM/E0lwRhRVwb/E+YAQfI9uVzHb
bf7IlE77bSA7ed0KZW/LiW/8Rz1aA8OMSHT53LbNS0sThyxpF5TdQZkDI495ipNXKjf+lgYKAOTw
Gv0ok+arS9GQ6/Dp8FvT8/mCHaqDrl4iWrBxsGbxZP28nCkcEcpzdtmytexWu/8fr1TNDauvQUdQ
YNnFxGZkIXuRV+wseelj9hpicaIkG88DCA21+6VM2NLdfASnkMUPmbE6bP4ssQoJVk7yS101qFUS
FOLD2f2qvuid1guq4yfnF8dgoof1FlvT6tEoVNoncFAh+WB8Pbt/MZIFG7fzWJrjvoTHhLwVEBrz
f+sOgQvwPenxCMCtAutI1fV2LqQw1+USXKRufrqVhoj/SSSPmVelFJE1pCfeEVQiqGLZDn/pP7/g
NgNw8zcHUIYPf9NDRF1UG3S0hjJC+3BXYp6Ck7955mQV/q2s1FU+JWKNiI8kkx8I1+TNoxljUqg+
OxPKzXNMSk9mtW4joXROliXsUw7A6R56tM2UoLzS8qeFVeOF1Hlwsblvke11HrRMJBUDbyUhrtPn
/EVHrXE3qbKuHG4IYO+IQ5JmXRQ5c68hgC7m4QJfhYr3LaNHo7OftH6JB8FPoM/rcRaBvJBAmRLR
iniSNxi8GPCYDC1EFinNyzUWNGPIFdC7WxnVMvn+V9qEneVRZfiubCF9S+FwQD74rBk+B8vhi0xL
3lTTarrB0SOVjer1F4f2E5tO9KBnMkMxkoAH89i4lD/gTDwG3N2iPTMkOcnSB7rCOod/MMxJsVhm
ISy1Ub2enax/AHXGA9hSRodbHDjy2epSI1CjUnGLHioCFvoEnqgM2dsOj6Pt27fwdKjt0d4xRCHC
dmndyPMzrcmNwq0VypOoLqfdJlR8C1jJww8pS/3nAeDSkqSAuVP13+3apQLM0Hu+Mv5pZpqXWv47
Ce3qMEQjwb1IoCw5rgsWOICMIhBArsXPmjoiiQCOadr5Zf96Ghp3Ea5CEd4vuPU4PfCkvBVNDPsA
KU6I+3git5Frg1YvZWNdZ9JQnRk3mwisRke13hR82pTW2UyCI51Gpz1b8rnAH/ukpb6c4zP8G3fp
p2LV474lAlJQ+AxFKqF6xwwUGYUN67q4Dly9EYtrJnZeOTmImDEiJiCKxw4XqhqVWHxA+/Ja7byj
1r6NTGyV5uxaCRlAa5C7wiPMK3MkFoE9knKUbxyZY29XMhFnPcZgVsAgRlOQb6GWula1tIffIGdt
NOd2XDBpu3ZMmC4mnqzC5s1RkmUzWQqZzXaI65qGuzF2/0b1iqSFQ7HCn2YbUH94mTOHS5f/sDdD
8lw+xV4dj1dJvrif5qmoJw5upQC8nPjJZkRRcpJQUW7ky/738pMf5mD/m3Z8ojcIqTjawejYy939
TDYl+AaE+yZOfkeLvHiUEafarcn7FS5eoBFMZBbheK4nJ3t1SAsH00P3PGtPxkC+tAkMbJKRUd/y
LZANJ1Ozc1MBoVIF+FRIIyAdRv+NdzRWAT9oCwSnPHFxbwiVturRQZ7tMfrlkrV9rBjTYqNynd4U
CPFMjtz6A6t4VUjuNqn3xdn6AHm2vAYeuuAvSyCpEKb34MyM8H/GKfTMea1lCVMP11Buav3qeyk+
18l8wzZ5jBnoRaSxRUt5WLNRHQUOZ99Ng2lBSDaXGGntY3VphjzT8gPNhtcb8VIGf3kI+MfIK9ny
d2XyOQ553Ih2dQOb1/13Dw4lpmLr7smPBykNHigbztkPMGGzjLNcYxLg1Bz/my5xXIFoJ1GpRWvm
JUel4dTFTljTLY9wiaX8tEJSSdrerNPib1iHDKiq1e0ls5ckVV2Z/LRdR5O/mBn4776SUw03NNkA
cHWxCovQ3dTMH5Sddj3rfWuBelRYx9BCHhQmoytYj24Y3InGg4bms9Qpc8k2XZlIvbV+hZl4DH2i
brL79rftN7JfD0jGZCIjFVAng1j6Ob/O1SQQaiz2SCMzTPYK/DJHrm/YKuTvXaGZLS0dRkEC+W6i
Nu21+DIqNazjyAxkFERJLDepet/3GhthfCBxr+VvGQP4Vt7Fx8+IhWGbZDn/OPZAVkgjMaJd3nLr
C+aPcpTrmrrba94UeqN3lYD5/qfljl8/4+kgnYEti7qNCrl7XWsBl6gx2c920ECesyrQuUB39ZmC
6uWTwQSwAoFmLfQr8yJKVJzuOxiazu5KLxgwiOnSq5sbwAIGju0pRihkBF+ljjiYv6c/dVKSFkd+
1sIfVjilBYCBkiTEur7hEybCD/Ufh1BZwmo2iB3TeKSZcresN7dHE90V6DgVsZBLM1EXW6uRpcPJ
gn/cxAy+Mamo22Khg/+JSVxuap7ptSu/YUGQQJJ+j2X2lZOsBjPP6SI6j4N8RgG3iAeM6+lrnUVU
PozjagWrSvQ+IyBkNjVWxe5sF/tjtNb0K4VksvwGJuiu3SVCCG3gTnWlsteZvYyJDhPlQt77uh2r
vefPBWsmETt/FGcOmJu+CZUuSUy4jLfVJrlnSzZ0HCUZu5dnbvgcejOPv05aKGoBXe5Hwfjrfcix
JL0YC6O481RiWasQGc7VXTN+/ac1+qaQDM/G9yNHqGCn6Oagset2URRxZdE8k0DGH6MBL1lcBvVE
fefOtsO9ucUokekd5RRWu5026QIIJ72IB39X8NoZlxP3oSlRq08Pz7Oz57SWTwY6FGxQFHprK9Nh
UilLklSXs7uShEYKyaRPC0ZVnQ8d4YM7mDV+ccR/xqw2IHWl7sqlM0O/flkBzoNCrVKmlGzl10t3
zUk38wUCW3QUPEWCia/53sCTQJdZjYOhDgIPLUW0pZ5yv2lzcFReRjfL9mEUdIGEcvqyVy80B9Vr
ytEWiJzuhUmvnnvczfwlZ7XDeg/wzOB+wKOU4pwLLEsHhfbAywG6RiUFM5kSYksqeADww7mVR67E
PX/xFp3bKuEpSsTdpppvykD6azF5pzLWM2XKBnc2hiuUbL41Qqd2QlGtk0xHWKFa9pUiWig99QSv
wDyIUElwPdMgJAJSlH6sWFTXBDIsco8KtN0r4RtSdtTvCxjbGRVeUrsjdcvBMSSVqLGv5VQ64l6Y
M0a6kADHNN20HfC7iDWFGKEw8w9Usze7aQ2Vfjn1ovxtKUAk/WmaK6hJ76fHzDrHWHl8qJSzJ1A8
0TJpHAVWiOsgFjTpPbi+t0NIhe951B+Ue47aHDY2xofYhFwwV3QsFLt59vQLpud+WBolLhM8L4KC
C4sPYS8GMqkR6lSf14gOj5rPvOd+sVzkcrvCzVBY7vIPZSjtX13OizILH6Ks1WQQB4Tl//xKYyYj
yblJMEjO2QUdB/CW19ON39owpt9c5aY4eus5Ri4iRrZyrFMwbyvmtyP8sdCC44XzYUppT6poAKQe
ryGFkSbsO6YheRayBGohhkS0oV+qyoeEWQgNJz5JMhsVUrsxkl2olHtm/OfN6q4tF37C9U3hTZnP
CpE1R4KMlqh4o9rZQT9PiKvZLlDCseBnRcnmpf31CsJ7aT9RvvwkqQlOAKweQ6yw8DkL88dUWlR+
hkGXse5udMGomrqSul1Zf/RY+pQyH6u8LjD0pDSbEsVIxx+wEZjWTOARV6Ydy+iLCxGfEU3Wu6DW
PpfpxXTbZl+6I1kZOUnh19BDVIiubHGqZxsXn7cLEiCF78TLxRhSWlMdZk7loGyxDOo1Xi92XlBZ
RnzoSzZDuwu1w0y6mGPiyFPATiNmpPTWZ6qG3DzuwUeHKrXkL3whgFERLmqsSr5nI6LjqPtdXxop
Co9cHL2Sk2njg85EnAJfxu3OTuto3Vy4Ve6nimdm+J6hHONZ7zDhl3cqAvSFGCcl4Ubl4Xobdbz2
lLxFVghViWMh00VSpUshtPREsLD5cmjmF3KIjBU1Tr4ogHDL4ALHc/eRuFqdEfWcdo1pDkDVzOxL
F/RIlCCiay9e+WEzG56iwqXbedO0jIZZvKI8t/CyMr3fmamJH/38KNeoZON+AxX/jknAXcMoZOov
7sBLcrQcrINb6dP4CoqQEOyKJBy3XiHbdvMqSfp6lBJYDlJuMadWKdMjXWB0Z2zxH3mqap8KUFWP
QvCYiueA/MIniqhCU8zZsA7yK0CJigvzwdZJ8SkQviT6lpRLrI6vYU1M90PYBVaAkwc3pmdx+Cuu
txDwF4OeqH6I0IPghrTZ8/TuSTsjfQ+oQ10r7LEbkkXP4n7kmMUARkn6mSmjgpNtH1rJ3GkGnqs4
yqibo3kdVGELN0+3NoXgBSPSu0FX7RclJ/EjAnkFHN0Cy9ZAv3CV8VgaJ32/nuV6XCU81XYdzhBX
S3FObdiq3LUBV0eaFBo0DBqhwrUonS/l+J/6XW+z7b5ABOgbQBZffPyxHoFiqrBdGjP563ApFb6p
5g43VkhPK/8wvxD9Flyqi5PToaZpvLz011+KBvTWyQwZUI3Jkp4aRO7v4elwzf/CQm921hxB1s8k
si0n/ci3KEhoEdaIq5rs2JZc/xyNzau1ZX719Imj3To2yE8Tw6br+QLTeCIQH2mIUFu1poYOqiuj
hHuTkrtLrkHHauUnGc+6UKEcZgx/b5CJOPfKZ4CqDaFxXcYDj7bZv7rRVoMt017sZWtmYvAQ0POD
pJmPlkU3vFaEpXjuc9fO40l39efAClhzPbOA02iJqPP86TsldjJwx4UbG1TTooK4BXtRHrwdbD9c
ibIe4wok9kIdqi8A2nmT63YVJuncAoHvBiv511szQnXqvrAqYHqqlZPsleyMULTNfOwZ/8d3ZnO0
u4aJ5Sp1/8iSJf1hT2QVErbsaMXHAR8PneEwIkpS/5aWg9RyR6197PZEZATp+I84+4fgsm1SAfR+
eLNI6vM4Lsq8DDs0AZmRrwa+h8KW0PaIP0+JewF+ClIFnSyoFV/wropOBPNfamjocgpTwCUCRZ9C
EAGTozagxNbsQrSQb6lc+tcLJBu/t6VY9kdLuZzrotsLaVU5CBfKEkZjgMAORtQYjY9rDvIVq+gC
GZedRCuB4bsXC/2HuICaJJyAIrAi2+PZAKudw2VeuRUAQjo2ThqFME77al3KDT96EwnLzKs9ylPc
kCS5tYbH0HkZ+BralNJxBO9n7CnILgWbaql0EKDWO6aO7hJ9sQiB+hKZ48t0JX5va81IwceZD8Ux
De3vaiSqLWUmGAUi9XlK9gPk9DLGaEUZ7cnITjBjgZ+KPu8xKWqcc6ftjpSNNE1YpWAMBTdGsFhA
klG0/u0skOoy7G1F9WxeQxLkBGjzrToHvEYvJVuZZOodyklSolxJvtCw+lwr+TQCJyrzuOcwUlPL
QrVGXI1GfgLa4vgucxXXWT3T/RkaC6L5SQtCNGdv8s8EQqj1tToB+cJwNkeQpcykqc9MGTBn/Xqf
nsYiB+xfpjpJYfxR3E47m/fkvmG7t9tjPaTKK8189Qlsp8XmUMKLbWTxYYO/yD2dp9AaEx1d3OkL
3QgHqKfcoPU+ncjeoDi/P1wx4g+3FR71IWA74z5LDWsUGwvLlu6yDcTsyjhxVOweLQZRH871Hxfh
kMPXEOR4VWnTaCFRhSPFQS3OXmX22q6Roo1/j2P3XmDxjM2qwvZ0ENXkpewGeoAtCqvwYjxk8VLw
rMABjpq7tUYycbJaUd6lmOnG20YZl9i5NguRvwHxxtMipEqB1lohjM2oeH36W1ckVurbUESIoPy3
GcapAt/rtpsEnwmC2UPKcH4dGWLYANlD6zl0aam52Np7pOLEbwXCv9Nn5+av71X9hF7exIMIIzNR
uCuR6o/ErRLzD7NYLxmkGWai0B1403zB7tj8sBUSRTMNairmyN4eboT4q2QWDAAiXj1DxbJv9KnN
sl1+Mrz/D33cGrZ6w9u1w9C5cEPj4ySNut6L/Ddc79zynF7NUZappf/gK9aZuxYkHVkA9FJFd5rO
D7LfUFr9nJ68JbvHZg++TazN7WfzTd/ggcs5OSwlbwFsIoLbQq8l8AE9sNWYJux2pJ5jMAs4P2EI
MuS0Z+ETGJZBtP+Sn35C7nL8XQ+cPFCIKdjAr8mbU6uzGMwu3Yrk5pDtxgd+N2WcLY6Jdv8RHx5x
+GexCel01t/cnRlq1Eed+WtR+GrcOEiI3Qv/Hws9oIIj5QC4vbrBtMY673zwLmHz6DqeCmo6H+gt
WRevP92I7ajc8RVVhqngxAtw1GVnJCTnFXLa8Mxb8ovtecA/QZDXo7hftDmXDma3y+m0ivl2F1vA
j3V37F/6G/yo+pQ5gVUKLmTWPBrylYgDxtG0+hzwLPz1yWyg5chVGW6At7GxqSU7ueuqrbU97UUv
HVYwpjeQgUDYsdV1SppTd/iB+yWaATs/cIJTAZUIsQhFzS6L8aCPGV3EJ11Na5pCgC1jCy3Cfizx
RVuahZ+7SvTQFqzLTjYB5MtgfGK3/1MMe5kPDlpxipqKx7Q7VMGUuszzo8QNszefRnZn3YjzXlDp
zLww9xaZRyvh9SJrdQC+0fnIQer3cNlWZbc+xNHw1TFWq1bGCgoB/nV4A7uGm7Di3qWaqGpfr0DS
kmhVLBftujtt8lQ4d8+X+1uJOVc6hzGJABBz8sKqootO0CZmcz9AzOMlywXFLYZ9AP4e5sjtB5DT
MG4gnl+8uVhYCW0f2i2emqCKkOrLbSfyF5cbbCh5CAw90qKyfeRjJtIkFo0QjfbahWwHZ/3Blm63
kvsyKt7isLrUVJd7uclwjjwoS5A+GeIJO1BlVRX2BJg13dk6/jrAOPM+HEK67/1yfB0KFNyLAQWy
EeLZh7/tGgrsu1y4/YXjwMUSiRT3Tn7jd/N+U5SiryDeDk0EppTP1+4yLV9+3oYuKMaRvkNSBIkM
ylLigjyTTygwVdI2v8kx+Gt3r+NbM22ARBN8QY6aX006pqFa/srVei6kNQi9tlgGc/jyfxtIPSKF
Ie0ckU6SB3R66vVKHfJeVRxTh6YvnLuf71hhXteZbXz/Hj4EzEwqmr8RnPDKdXN5ckL6ugDHtwsP
cfNz0pXkP2QDPUr0HOhjddKpjzIY5JFNoQItEDAuW2+K8PPJiHu40oo0m+aodd1nEMhWz3uHUD2g
4Vcl4wFR5lYwV4Ao0qcjmgrawweuJZOCbRL5POkk5LqcLcPTVlbd273auOn0n4y/v3ix5yJ1BZdE
De3GN8rOFShdybN+pDhi6JYAEuQizJXXjGHEFAJI83CHFPlrxIvCQ9QbbHiKXd9iBkxwOPrfR8Bd
55IJ17FnuyZz0OlIBmT4at3fb/IBhPz4U8DwkOFLLHlobLnX5Y1a5GdegJvoa/TmbEjssh0ow/+f
Mr66xEC38sI5uXAhrDMwMVpNGl5EwwK0Fg12XyzwgahVSHiAy5V+yadmi3YOeL0ng1RNbohvEvnb
qHxlJWvGjmWTvyLHZlwNIYAnnpFQD853/ydlJaLfL9ey6PFEMjBGBI1ajXg83ikc7fcxm7mcFr56
zQtdF/HsiUTcZHiV+knR2I9ARzSgE3la+8FFPlUy/H3QdsNiGG5J8MoSegZtqpvsIQyg7X0F2rmg
LuC72QEqd/SDZdW2H2cwAaA5gjitGgTlo5yIACPoIufLxGJOy7f6CDp3UaXrPqJziAS3UN3Dmzr+
PzDXJe/+wztzuJ2vPdhMWBup1U/Lft4Bzs5AcDXZb2p6dw1rHTEzIkOkk4PM8+NS0m5HwKsyFvZX
DrB6H9Ha+6H/ZHIP9rjg/n269lB2x8tX+nOJIDvWucKq6ZR8OQOVNkLxoQxccx8VjeysUKAaTtHN
OJOpg+noJs+pZv3ByrUvPkEs8lnQZHOV0yMPlcSkeqPLOBROPZbumhNA6oCtzykvEs/RcLs51Ubb
RgQfAhLzkJCrLpD6ytLeGj9PbrSgFQM5TeiEohvaaaxHg9kbZgE9gMB/G6hy9so1Py41QxoobPrh
8vqyOF1PY5VcFNnBgWcXvd2V5hvbqh69cW/+cmaZfepJvx71srLLwK4snuf2kY6mrMEkFjhWRWwi
vKgT7OIs8bvkxIxviOwOzZJXXYP5LWeFJwWyLD/fmoWBoxgRt+eS/3XQ8io1MRjOgDZo4pM/elF2
R7uHGe/8gysdXJs/7J9rHuTdL/sV98+VQaYOGEVL3e/GvWIItsI1g/WzhAggJ3nheTDtF3wWOtOK
KVB5udzQc57Y+XEEAgVJywJjDZOh7bSkTvB9/KyQY+ZCJBKjT9Dp8ZjKi1EJb51VDQG+Q1Y523oS
59bnPtVA+4iJH8FIDLmCQ38pJ6x5rbFgNCq2OJfrY6cJ3pvYGq8hOzpHaz2BmU2YKam74gl0gePv
rMymHu6t0pbev3ONj9/3Bq8h4W5OJDJcuiwZntXlkjnHwBa5JI5BLbUUh7x6E+WAooUt4XmnaJBJ
rN/520lR27DbjPhPNbHVsuNvnUSSIKSSoGhwVRErQTNgiad3oBg91ZlielMkyglyAOFbIg9bJH0j
QJ0Oq2mQIUhEsWhHdiapHFsgwKsOkxxb4k4xdBu2615/7zWIV9p+EQOuwkt6mBjEHt3gjvsvTfkR
k9GOJjSHk4e7IDX4XhcGEXs+TDR1wtl209pyH8XIwS/CghGHiqUT2ldHtvaJjGqsiM/5kWPMDRg0
FVtO9v83gBIxcMB6HShy1ZRy4WjOz8wdzk7fh3wzuu0Wjlr6RnZPMBqzXoyXNUnVqrQpHgxi6/ge
tc/2xyThO8B59Kb/vkK6NEveZzEEq/WQLHAu99IB3Wc9UASd7txh0g46IXz1aV4rK6KxOTbISvmH
r628Rkw59sXZSUssYPJ32StsILGKNOFicgRPKzoyfUI3prCyDmyQUYS04twebaebE1kmf7Nq2Uy+
nQz1RO3lAC2TWXRjY/6oz1ljDxwLOtlwH4EWrFZVu8qEGgd+J2Esl/5xW/fdrmhrtr7/L1kfbnyh
pFfFv8SpnwJyoQ/xkbtmUPbuFlGvsHZU45PAUflxtyALJKp7SCU6DY9aIgMfkBrPGxolWlu5HzcR
6Sx7P8CKK5/A7Z3Lh1Hj3qtLpXYy0pNaQ84t3UmwfUCBIWLtldZfepAjeT2NyCXnV8DcwDgfRa7J
IRb9hUQGCMExof80220r5aD7vSVebH3sCv1Gvw3AX7eXuIZtsCbmvUIxu/jC/+52tSKX21JHFNeb
PC55mIZw2B28r9/1I0IDWn7NbmpiSH0tOL5MdhbspiPtm7vjAGCpbUx20lejrSDayZsNq6LTRjLI
5Chk9iGYN71qV7qmFiU7idDZOz/PwWYHR2pjGUS103hDZgUc5FqHnjP6kvonPaJSQ4qagJFXS7g3
JMgojVEf4VPseyWpFnjitQG6V/7z0m0wSZ5yLCuE5bxknJuKKjrt3MMnlP8Q9/FUNEuzfhThv5Gf
Xs9Xlje8R1b4ekPyKmB4peW+3fVs8QwPM++ogZv7x9jGxPVe9jrcQjWLn8QWmGZPjeRLOsgTCP4/
PPIAEQOAQ/lNRIvdC5hWTd6p3KbxAHztky0UiN+UlGD8+1NRvqGnL6AbChkDNfCAvOHNXYvrXz0K
VT0oDYv5FS0V0N6GkLLUy9UgFbKekdJVRni9sJopDnZrwm3gKSY8366gbBLf0UsplNVlNA4rmBY8
I9Ug0iC35M6lXlr00l7mWj7VgPE6Gqmzf8SsoKAudYg9KZHt2PnjXbz5JjlrrbvLQhyoqHGV5lvK
0ohC08pjQw9U//HMQl1etyfC1elYMqtyoieiipBPoxQRX/e18g1ZLRPZIMvR0oQASWKHqicVZGYT
G+U3RN5Daz02K1GE66amwaaxSa5ujzpAoAy250GxCdgWYlP/RE8wfobJC9o1qUbvLWjXJ2Qh0rOw
ZmXhlV8pLrg0aLkOHjKYvwHUKlXjulihDtocZYF2d5BsP/aKylsGS+5fqtwvBzjJRwsDVVwZacLc
huA+DoEpyJ5iyKsvZx/PzNSbcA15aYdQNNpkUbyJM/Lu5NhsTQu1UWAqMW7i3F6mKB4wb8aVpMrd
w+O0Kkd6xB04gy6UF2xGhYyidffdZ+M06GY+DemviKasYspinISyI28UvGzyW74VBQ8jXrhUL8tO
TuMMrVPQcj7Rp4nQMrL0G492cJxJh68+qvxiMeqH6Lfd2d4/N+WDdI3sK/zBEi0Fq+NqExI9QovA
CsMBx0gwQtszF3J668Sdkewd3suvrOaQcxd3l6MMysGf8ebwh7w4is/7TUzS19VB/k6azppZB9ey
GrQH7R/UV4CvPsWWjusz0HZe7mp7ZnwoeD/YQd5yHLU8YybMbfKtSMuJW0I+rw15apdyigErsYBL
nIvUrJ+Y843y42TE4akFDG5Y2U/H5foY/T1Unt3oYY8oZWksvcyhU9sehlhh1mvEa4RwhgcNxngI
ajzhFIl22woWo0FibDx4KJJ6brzI8eJvOH6uRHbpQXfZ+SIItoIkK2ObeVA9iWE5/qaRIflH6EIl
2GxxcMw/nvQcUEmyKx73tGIGDQsdomtG42+gE1M/CEkKOEmo0wSiD7tjhVe+LG4hFE0Pc3m5QXUc
v4hb7cNIBqjxyaeneoFoS6bNB0d/622f2EKPWSon5WKgD27MFpIX//iMpTgh3xEKerkag40rzrW4
TRmVC4AGxzp0lF2Y17Gh/HfPxg6a7+2ud8/RrYT08bZBlKHcBjmwfACw8MVl80mhn5ZfK9CUaI4m
b33tDtL71uQ0z6YAan+oKjtRFDJdb4A5M0hk8Woh0b3gsHoJIvZtaJJJwOIbKZizokU5VNTSFJYW
qmFPd2eNO2Y2SILPYU0U2mkyVvc6g27SewFDTCJSURa9rYhOQ15tNv9WkZZo8OjeWSNXuVfTFS9h
eoc73+TZh3iByb6gC3Klt84nL/JX3shBdbrxVSZegtbpKCqOM1XnSTDWkVuD+nuRkKGZJ+d04eh0
3LYohjccVeUImR9niyVvxm+cdIHuxNmtfx9OYDY/mlK347ihvKOvH9HUT7VCqKGoETR8WORpnH1f
SUUVl4mL7QXbbOoG4BafwvT2MWKpVlqhkp9zI0ocZ9t6FQCwJBz6UDTSXDUk69bKekN4GjgOxdKm
SOIrlZl25YTyCocaBC7a+CbtgFV6KeJPYfXZ/XYbAYtEOhJi3JaSYJHd30Av3Q7HGw5t3SZeAhee
4s6RsxIJUm3RIRT5khcqzEzVmhj6H5F9fHYnBvUC/xP/v6wEm+2ZB7qTOMP8s1PjlIpwhcFOHlY/
iTXt5enBbTOZfkQKr060sSZIOKZeORZATvUDpgKolRgnJfFZAIOsj80qpO4rQb1dKFivDZO7Ztj7
fASROXQ7uKOFFQcS6fmhqPomhgX0PiwolqYDo+5fiMTPT5JwgSyDPbSXbBIyQHEUQ0wMzItFV7OW
DPwK/tFUNE9ypgS6bDOcE2hDf8XKjQDfsiB0x+ZngffHT+y3X6IQ59tQPwRKFoKYHru9SxI2wlIv
aPDWc9or9pVQrRCecUh2rVbbWhaBAENJd2lLQoo7am8kaUdHlrplxvT5lPFnPvPvddkWdA2HZlXG
yEZSKeBbkTY/l1DaxqMMG6HNQDYIdQaq5eoAa0MTIcK4P6+4nRRYQMnhSnlkBeHt5lqIMbWIk0H4
Bwxou7PbMUqOhS+PDZULWtY4gCd871Bkvr1eP2hyVAokB1wu27J4Fm4dPObdd6RomIJM715NkjAx
GeW1limosrU6H/DApMXfKQSPN/zDrb2qkcYJRPIUXaq1+h4wgbS0H1FChIPPIonXiBoKdV9IVZPO
aZg+p5cOoJJiIzDWCFn+odAF7+2pdYFMuMeFIXgxQ/yEE+sAU5R4j7EHWV+UAPlaeAErqPIb6qJA
mo8oGtfagWaFPCcvx+h07jMmnVF4YV6eulL793IPaMxySFRdSzZjGveXHlod+kkSEDxP3ZFtmJbn
WK0FTiTjtTxvFAa21RaJ4fXPwN1mo34lstCIeRnibfY9ClByuuP7J/ZyMjjYuBChxPk3HWAkQ4tZ
PTGMSPrAvUNDfv6ecj9VEYtTLtHckA9/CMitTPgNVZgInG6Jm+9vFkaSgTBJIfjWO1YSs/ebUpum
ttqml3/oNMtQj25S5B4F6CRTEidLv12a8KdIYkWk4aYoNwFXkOSOwQcE+Zrz6+GnDJqULG7so3Du
cj5+PVbRF49vCKNAwIMv2Me3bqeCCRiwkaZoJ/DQ77vGGSC0rIxrO172Ga/5Yw1tZMmycAAenbvj
ttQase1w51dn2Bs1sa83Ir5XSOXoV4PtoQLLC50K7taJJ7DXfdvp91P5T13oxL5miI85rripZiA1
XjXcXrZvtroKLbRsk3Zl141QVtHk0el4LmOXG40yhpSMa7/DJpo55z47dPtbZxG8cPBbP7SXkM6Q
z+8JoYamswzV3YWrSoBbnp+bLQiFyrW/ue5Qmsnk5J7ssu8oBZe2rKU5Iyuu4ezXVXS8D2wpS+U7
4K7DRC0ALCVLDSRhvTM0WOgX6CaeewEIscmGGD7SNlTYeDhtdUiJln9ZnIlpMnUkDob4BbwYUF7V
l7TdsAd3jeNef05Se54251UZMFS+qSgbhFwmG6a7GRiNYzxofNd7BryRb8gRkMW+WWjQQAFs8FtM
l6YoSiMKNN5pY9ouXFQW3/+lP6iCYkZ1Qn1vvcXZrWDSUXdvRgXicGsLSqpOD9cv+kAo4HkPtVVn
i19mSTkZwbMO5uOlj7kwxaQUkSouGwjQrWgooz5wDcZH9JMjo/01xGQrEZONKghnMVpSAVSWfWOS
/KKt7uklmJHel1Mvmlud3RIaFUAKUvN6ZwC1vMB3ORAkiwG0rOGdfNZqHboCui4H/W8D++VU0kRj
9euXYDI5VGsDbMncmxfztTXxBk02ta+vn4zdRZQmHM72NAuA7WDX8f1gn3aI6qCdugUji82kWV3N
2rHswnn0tJYNhLlrdIRyhCS3ASLHc8cbfbFlW6MFOWqj3H+U3XHXSfnt1XDhJ7ywe2yBokTg6/kF
SBF/jrEqEG7ZL///zuui/vBwBH82WNcM2CKvpQWu6I84fDMmusxP0+4x8aFMCWlt6WViKmCaCPs2
DRyOiOUNvrcSCQcX+N1BmEvMXXgTJ3BCy2ruG/DhE03MUYhSHjjgiYdlDayid6UwfvdUaxvp5emu
d17CvInmE6BYr6OR4cWaueXEJroUbIcC7xQMq237Iw1+8kw1wr0sQh0CKeb39St3mLXQt67bETvm
LHrlSak/c8h5LoUBGNEUiixcKIfrLjUPmGc3VTHGBWgRdkFqREfoT+VVM8X/gAJRU+UvVea05VSs
W/d+jgTBtEqJeSffgsG+OODGzfR4E+3C3OhiRc/PR3TRmLKwfQWoRQC/SFzgSjRZPdtTsjW3fj1N
reSmz76KK5fh5BaYRbjMyJBP7L6fupwWQ1tiva5348YcgQVVrpvsCpg1E2pqvkYj52BvWuSxH10D
EkiKoLuQoS+/RycggQadL9cIcT6fhqnjB9vDbu93MlZzjZe+6YbdX9ZapKtdQFHe9xKvVNGdRZQq
pnjUwOhUluWqioMArqHCaEsHXQQSwJvo9OctmoDbTzu833JegvPDCD3OWGOkQ4YRe0G6Nn1GIb3w
+y+LjvBtglI4BIilW2Lhi4F8xc47y+PlJzKVuGaPi449xk4GIbMKmTczIIbErZb4aK+Oyrd0Svn0
ne46dLy14Cs3LqWpp9k9mch07Fvn2aVMyfGCHH8BZ/drCc6uz4cbIEBA2N1KUkRkwtYNYnChSKz+
+nzcYyE63y+gNwOB7zIB0Zcko98PceQL/CfyAXcS3neue+TPsDXnUTZlfl8Ck5/Ti2TB7rxCp7au
SACEFm8CwPBzt2sezgpzzA3Jk2D3/p1Qurj8azP2+q0XwRUYES19B5vRlfA9x4g7BCUxIgcLALVi
8fyvrK2l0kyuIP5gZVPh7n/aD/wyzQ6GTjXUAyEBXCNi4+mxLjBcXGf6SZWcT1G5sblVb8OXAIR1
wmb6yerFO6qxyUJM0HUs2Py4kS6j3j6ZsXAouVffdL8HgQjwEIPZyiOV6wg06uQye+YQ4wIs75IJ
wVGa9a31SrdvqlAFJGceLOZG0iXsn5RYpUBGs4CcOLEG/EG9h4I7TEeDAG6TJWJLuEQiaSjNqps4
q3sAtM8vyB6ew3dN5fhni7qiiEaiT0WPGdpr5vVesh9iZtjQLrW/e/7rQNH6ZlFUgIJWRYju2Uvm
wzyTEaH4Bo5p42/Z/fQ7eVY9y/Fl65RUei8rXsUTJConJUsWO2PKXz81R/2G2yc0McGtu9RPVYQP
3gBIODzla2Js611AcXABiwdRBwfLMS5WMx9iFw1uYVstyA4nykdm8h29FHg9lyvw966cibSqqzTx
Fl6aV8Bdelrzx1d1eUM0r5+HgFkho79vqLiSpjbpCeUZTFSsg3+ueMtjczQJOir7AbNVgQ2TF3Pe
S/EjskwAQDkEZOMT/5KTFnQjQFoxWc8ekr8u4//wXoivW6pbRcmYb+NXlT1NSjll2Ook/4mFErMt
03QBev15a1Wo5v7bFAGN0zCRb0u7ow1O5yXzSjDV3ngCJ2oWhMnNOYcTDZX2xRhUs+Zzy5nAjLda
XEcUPhAFyPBdaRjpcnWyEXlZUsJUAKgc4blYC/hgvxYKV8Jwy8xlY8jPvM3MPGpxJQL5MyWbk8Zu
RBwaUYhlB7j/NFjmwz5uGgG0c5A/97hES7mBOn+BWST25DWMrjqhBQZfmsFggSgMnnJifQZEOMJO
sB05aLmKzxS0GwV+bij5mm6zjenOScMjQdsuTxS4kC6eYtTh8vt4hSlDWHqwgSgXzEhSOdLqiEoR
7sCdm0y2j62DVVa0A5QFc0Ggu11mef8mLOmL7uq5nAKP6FADwHkBBas0PdKblPU6HSBAFPJdZDEX
dE/PyeZUkcolZfweVt2Mwn6Ci2GJsI6FAPnUWjkGqDMnISUI4fTKZLHiecl73Bfn1mi/wZThklRa
EifAVzHm33IcNCWc+evvtaRldopHlIcqd43fQ12tMmX1WdNEc3aLgs8fAQT1rSDAWfHb+C3Mnsey
0oNuxB2f/P/uaXUgM2/dVQro+mA0VegvJ4izyMNapL183y2aD0wYxD4t/1R0ZYO1BiT6sGrgTlfn
gF81QsX43Rn9RnRlFzL3Rsdl7tI3iWRgRKzMwH+GC40wr5m8tlhVk5MwlC2D9jH218S2XiiMuOto
qItAvXdrzvi1PPhLXAk5RrcaFvUn83e43PuAXGp0oX6xwXQwmpKsK1J4vzPqv+gzRpyQgMSXeZgO
MGQORneF3WRE/E+cumuwOq6cUagTXuWrkgvwo86xuJlcVQCgHNAPO/z8K84p83eKDBzXqe71IaZ6
dkRs8SUvr20CVDkX00j8fBxyw3IrTgKe79w9vUFOneYsvn3FNl+AjlHmobu3Sr2n+iD0N2FoiGCO
7rDkQIkRlaVu02ITtqqJ5+uAKLV5UWLkriFUcXZbK2KITVnAbpbuX29g7VslYxQmE27oLBcDWetO
mXtdMMqaqBq07Ew6CObC3hHToF9bqucUWfvUECmMwiDhXuGg17SxMK97b12mxRELZQx2yOtGBpx5
CHeBqylzt5gRB+uZuuxC3tstR1y1qpToY/1IjO6OldAZ1C9l9w5ar5Z7TtMZC+5Qjde/zHz0wOwj
ul6/EAOp/FRidl5ktGJQeacopfT3oUds3IxYWa+ivsbSjjagQk9UbGgNBr2lqsQV6uS2/eRNGOyj
7FiuM5cfqAhyt0fTKgHrjY7Is4do/DTbPycxGj5kAkAK+8Z9HS4/J9eZWIoX18CM5JfEd474+9NS
m+FNbWf0HXB3Npx8Rv1hKUHaM0P8YDuKETIUIwmOUFrxAIg+RlG42bYXo9vsJMGEynOLJIFSTX7P
qSrd3DY0napgIMkshDaEYBKmj1m9bckWV4koWKYhMpxnNiTbQZT5YHr7DjvhEGKa75djYFXrHTsI
Wm4vN5e66TK+vnGLxBnZCRxc5t5SebJMkS4g4fl680Vo2XuudEMWvz96M6OoioJ8xaLY814DmUAF
qd04ABEde4StvYoQgTVupp5Pp+xJOafB2vspX+SZwbrBLJ2DLZhwGfF/r+ublD6rmgr6KbZhLEg8
OCAcB0yrISAZjEbBHUdDUmTtq+kReJC5/wKXOcHU5/9xd55hTBoGJhipSfFj3QzXSoKXoMJOPFrS
i1qK8y0WJqKnHUYUz8PWVzJKUMi0PGV+r9t4bTbBYVJJ+EyXF4SZ7GvjTF4WW0d+Kg4crmwBLFT1
kNnFVMg6dWuHU6v2v+CYEL+OtGBTSuFq/oE5h9kmvi1usfpvoJKHFegXyWabWb+2IT6zdki+4dGv
oupgD+g2aaaKXYUzHfOP13z9tN+LSb+jcG4Fbik8YUNvDHXigZToXwtRL06dR4SJdi6RaavDmUHV
xbarnKpQ/D/XAiVguu8ZeinJidNNs4cjQ/JgNZw1M+QD9mJWFkQ4vOhNIi3YT5qdLx5xAe0Z1eAb
N/CVW4WZntow2K1xcXmehW9eznqcfJdSeIBfr0l04if0T7iGbAZatQeGzJ1Psn4XTbEpkOYRJJl+
rDY8gs36rBXHrRt5SLMNwOStpRelObLZCWWikiIovRz5HdcuKHhaY/pUZ7w7scuJUf4QA2cp445U
4Ein9acqLAD3qlbcH8LhrIUI6GRcEc7kBkFje6Tumu5/RoN+5mN5DTm6C/rzZB1yRaiqJIHJgl/w
VU5b+4nliL9D4hEnzJ+K2xDfY2sLvl0sNJUsxipltD/xVY9UKYPReHT4ufQgUatwaw7WKOwRar9D
i23HLzuiyLyDBtc5TjN0snQf8Txvvn8A97ajRakLoiAOGgITSa7g9xaTkSTTU7zYBZokDCIpVTyH
ttCCpQt0bMU//aTWh31tQYXRpdjT+lf78serdRzCSqHsxALwdpqNCMakf4/GnyFHnHsZeo1NGeK2
tiv7pxO+m35KooT2QY0vQZeE0HCWh90BJ81JhS/lKxc3cwgmL3Iv1m7VB1Jvh9ft8vysYeaDzmew
dqsOZAocWojCmntuh7dLWhUjM+X9zZKmKV2OguZZOvfo5lDMFJAiSkF4Z/YVLz2NM96nOLdEJJ/Y
41Do6JSkrdC7ZNsn1f/WLSNdn7xTbeJNOfoPh3V69vAv+uIG5XNu4VzQ/YxCN57xpwSFhMp+LPEz
GD+hf+cy2obevDMBgkSbhj+co3+sdOFtw+cZzf4/YvCHgnVI7btn+rYksTgPwcSpAw9DyTHzI32v
t0ng8J2HHv7NepBllaUDJMyA/velYrNJfxlLd1B73Bxt3Vook7dQ1Qh8z0/9UHaRB7+XE/x3hRwr
yw0X8XfAu/l5qynkeHL6II3ATyqRLZAeioWIT3ve16nHCZjnw5pioJMnTsp8phosHA/5N6bhuTXj
I9X7BnBGHTDV+jUQqh4+LMaoMonuSIu/lrkrdDwdDo0mR/pZ5L/sbMfYH4SkaPMhA1JuVDb097Fu
pPjsPWDvuANSwBDOrlrES7gOOiGSd0cCQYe4fdihbv1sNppWBrH6aryY1VfQlZMU+asSYBm5KFVC
DahOjgBtr0r+WEQkznB6GOPPlAB85crU35CUlR2/MbrX7RubVULseEyD6L7yvBbCIT9QmcOvK9AA
9mDk4SkZA5Gj9LJ71dE6h0100d84CvzTFXSRs1drhjDiW6oLoT+vhOeH5Mc+BwNVFyv0XkBu74CT
8UfUqgWM1Tz/uaTXVI0RWF5nvKQOs11uDfd85J/RTsbLawsaV0VcxfsT4xWbUzW0TJM2vH2apwb1
LXIhUFVHN1BoqLCASB7LoUvnOglFrolhIEk5r3z7l/GrCL0KqIFkgby0ZfpZuDi9m0sdv3pfPNZn
XzvSZ41JK//QqfSX3f1vu2ZUJJ3nQA4je2rHHmcfvoDVk2LNsv/zbvTn0sjKFW+DbqYQxARsyfVA
9fuZ1U/MF5R4vU9yeN5antHw1lU50YhM6LwmlVppC4kPmdzGvfr37ofHUuPBRMU/aa9Cmj/iq3HD
JhigP1esPSMVMDe4mbXp4KR2MAJyIcJz0aeFZ9PI/Z+EXIXOBbFJP7Yi1Nia7p2lHo+i5DEyXBTk
ErpHz9CWIqLH+X4R6/TeETUVJHIgYBADYRkvx6BxDRWVpTZ29L6llfIoNGdxXcd8Km3MFctA6gsR
c8HWUSB/GASuF4yIseboaWV0RKGVR2H/1C/yNQ0bNsr1ut1GOmbPEcUI0W5PZ4JLRSH/eSmRelXS
9H2sbECI1y2upJawZS7TtEFrLg/DWMz+4gT8PWgJuF5OwD6M6jhFz+SvE3SCATxldP9M6viIp8uN
wBJeg8XJuvUAEbgnenIc1+gIFfTbfVLqUD12jdd1TuwnNzgrWSCXnLkc9WQ0o6yRN5xrNRTChXB4
vS0t6WN8pJ5yvgdR5Ws7xd1IFkJVZXd1nZOsYraApmh5X4L7MtaeP8b+KFb9qW3EeR+tS6sO6Tw3
lVixxxRBEvrLaRBkJzy0ywfmTbqUHMX/XtHql+cndmh54nT7+u/PUIYt8D0xt9p2/mCvI3f0XEPr
6k1DZn+BULNRIeI5uygzEMpYDAvh4QcGHLVSTdKxqAmp6oEkdGxlEnOpd6p6y2AfCzuLrFPxv3Za
UoxOSFkWdx7vHpFYrXXAq1xkTlJN7dU5SUJkYNudlQl2zro4TGO550t3PnsjA0Cl5b2jytKfgBjV
5bFDJB7YvdqtbOmYEdZVQYtruwMb7xdUI2jsNCTwydqlx39ADYEcH81ZsSXPyHxZiSNKV5I+A9p/
9pZ4dF14dlBN7Upl9KKLzloEOv9zLF0bE1f+75vBoOF3d9BRWTKV+Zr1VbIX+TVLzYRDjXhqjMC6
IBS9uOyAhWgxSiGVmoJgvyprA9F0Tcg38fMRuGb2ZVOCQXHoJve3LDUL+xTKB4s2QCHA0jq2NpLt
hPV3zMsn0IL5v2h8XOdsO065lK53EXUsM5tRJ8kc2xa0lFYBwn0IYdRU3QGNHvQaOCUDhmGWZRO1
erDgNJBG5K2ht+atMtemEcy5rbb3gtBvybKkClfQ7HF+lZeFO+enK2JA/j5fm4d+LsA7loefUCFr
CmpUrd79pwDxADtLbpAkcY515+ET+JnHuLa5XpOf56cgXLdQ8+qJEStDfR6/OLk7WwZS3OS2R2F7
QUwmGotXaW41cpWUBmlU7SF3K8YLV8Zgng4rRONORFDK9GTME/+hNwf6qxWGPM1ejIETaMn6+ZMG
orUABBt24RWbn7pT8/mnBOn/HwL54mGBK9WEorqkn9lgd6MvduRnblsYnydY0ZqxPNTM9v/gHBzj
OA95HuHc+Trr4GFWbNK2ycp9Ormv4/GZimwh3EeHtnfueRYQn1nCn511GpUBWF+AMp7ioqkD7jQS
qWbtFvnlsGqtL1k0ebYEOYrIYFLdrT51e0SB4jqRGrQd+HxOzbfnqjIaEh4OyYT/dURJ5qMSJPLb
Caf9dED62P2uYFKFYDhSIE9l3p8SaE7JbczKNaWAZo7nTxb1pyVjVu6Jo7NrzAnWopOoC6h2oVgB
kGl3WInOIH+q0qNCK0uWuh3D+i2Pd4V3vgMzqVl/jCzexL7rYddb0ku5l9ZXI+tb8QpzXES/OmlF
XNKjXUYzVJabGPosmv2Huoogcb+Ouxya2G9GHcrv0cEnhdp2x4Nju4c3a4VJB0FSusOUcpZMLUWu
Pv7qoMXS3a4YbFDiwZjqDFITyFgGj1CSbPaOKoNcQtrebd+wOOkYiGjCwJTnMIpu78+tprsbh0TX
Ac/rRzP/6CcCsweK73JZgg86pwkBOimbHAMjB18HuzSgGkRQ5esHSdg2d3NwV87gGeSn7HF9PviJ
PxjU3/triIwRLU5f41n6uomrrqv10rXET2nCKmKL8y0zW37voprqUWRbWKAK4UpP5StX3cE36ttr
Jm7LRs5naOEzdtOluJLg3bs9AcnYD/vYbykO5WC1F9NtpgoAG8TsjidkkaOojvyJ9sB4DXpWe4BR
TUT8epV/5H3w040Zc3zSN7MboE5ZHKB/wx+msT3UFDimOWCvS9d+omlsdoUtNIgxOFGvbqR2pfdi
KRSkfJrsruebRz1/6+BFTERyZlpRvCoLd0pH+61p6OafmfaMl14cGLJh2dTGqYR8o1mSgaHSogUE
XjKgwHFyJ14PnhNgD0CP8r9gLZ+2RNBvI8jo65QwKZaiz+xX5sCycJWYsMGW2IpF9uKAfQki2dn2
w3RTLkmyH4EVKCQVxKHSlf2cKrZjSBnSrHewVD9rMqid6rF5bU5Bea6r29qxMslCzDJ4+rsZV9ed
Oae4H21QjJbD4N/y1vN0IXLNQ09mTb4juOXPNi+bjpXKDNuVEMHxa9gXN5wWpxtexXAHph0eylya
qgXNXGukwD0DXw5cKvhDYaVvakbC4uvDlzMtI/m7vHPf+4gfBAbmt/FzCEm9lchnUYTPqcP6zqyo
nyzXSdKR+vKxUsp0bM+nnfRWs/aTSQDHWIbwylnEiCtkyAZnb8heYzvYuA7mK6xIRcBz65xvSgCG
InEBW/lnreWD3YqoUZKXEuM+HVeMpWFwRBURftneFuwV08J9UBqgFxMhtZYMkxYKYhwr4aagM1li
TPUn0l7BNBtJVM+Mnsf+qk24RA3DxoOZu1Uc/fflf//uv94ZOS7cPNmU/oqIQoi+YTIR1lCarcfT
3Cw40J01lHST0MHvb/8LZh7l282gPW/cdEADaGX2MLZJE+lTxXUajusmO5cqkALTASPMboMn0wOE
cy5ZlX08xa1obqDLHfOmLe1rZws4HkB0LhC7dHwmSlDBh/w6rN+IOnirCOX7qNL9X7QkEZnGe73i
Hlww/zkMSVa3lhY/NDpJR45ndbeIWL3RvuTryI6T9Ck554aqiH/7nwsJ1wxRIbra6vKfhfP8TQkL
gdXZv32mveZcTIYJsrmBhwNQbCB8Z1OsAVw/Zgi9a0k1THSbRMnWUpooWPiO+U9WSGw6Z7AiK6zM
3xAkUXC4XKnHTvjm4PtYTOgFJBr1ePRuTSbXwNWIIwE10aukmDhs9crRGCAnGJNB7XOWJ0abX+wu
oCMP1mDZBFKYQQKO88OecnXSli61qCqPKetuj/fcIfFo/pY8VkvEMy1ewP4aSSXeYvZChOs6GK1o
x2f6AvFwVGERaL8sB8aZ3nd8RSx1/VsMpPUSUJVSYGtgMkzg0Xxt9cVdalAIdpd1XEtFxi3aj+EZ
eVQJN/pM1c3djNSh3EJXf53lYfdQpyXpshTSwok2NA5Hi7FC8X4faSv8UtxgWBZlGdd1V0H1j7ke
cN6vg10TgxS6r3YLYqE2nwnj87keQpZskFcTOp0y0XspNes+o3Du7XfTRj3PRIfglWFkhmi70EPX
+jFRO0lZYigsI9yQrAKzCsgZ8Zx5i+tnN9skxys3+vfGfmxOEsuN3RjwbYrYEsFIMZmyQWK0IJBG
XWGxhH5xCCnJolgOdb3KWXjnhkLcv7SaM881Inz93PhhBQ9b2FFXuBImMdu8m4hH2XNAEvgrq5pj
rhd0Fy/rIrQipBoK95C6oIhDB0Gi7Wmbz8McfR82NlEgLdVJWX2y+n5uIWnbTg9pdX7aHEmbyIfa
36nCDFOx3w69zRtRsPEcDTVjA8xuouaMHiB1azGlEkzOB+nQGhsT/eAtElA48KtjlFqbKn6gNJcj
cFitnHPH+kL+vthV6UwSDBMdY+R28R9GObGsR1WIwg5YNEfSt8cqOzqQXoQU+MGf/eXMMQyO9IlA
MsiKyH9Bvb2agVY0E2Cunzn/xAjdVk14jjF3A2poBmXCKAzXQfeD6gypjzozuoMcM13GPskl1BjZ
WT7s8oTPJZdofZgp/SDME4823w5O+juPE1hDzIK6L04SrZapya9UKt+nnvszb0j2Jq9kJUriai2H
QiAu2cY/TCJG6+Q/Pm2JxkTtwRC8hbQ7D0r+GCr9YFsEmCkbwfk+Uq0FZ3ms1r+abNT6EOcHzVKi
aRS6aGDRSrWj5a+LpDCcgrgnY3aN/r2ep41D3o6UNkHlR5wuavPzKEMBTyJh2JBlaKOi9JC9pB8W
byRa8H0h2bZ7SaA/kmbjTA3EA0s9fw7+hlZ4QSvEO8/qbJeYhKqH941evwxfAW9DwExQAZQ0tbaD
k/ZRVQZbgLbQCpZ/bQqmmgnPYxX/UNvYxc5Q3VDoA2K/PIcmYf1a+oc6j8uD5qKha+nFL7RxnGEI
z7FCU8bDPkRFQ+ipsDMT/MgIvtg3qz/7vIZXRqHybg85fPTkuly/w/kmH+ymcb8Tgc/rxLF9ANjx
oMeMwpxp4qYy54WlzkLJpk2+p8Bi6+fqfkh/exHHG8upQs+UiyCZjSA1WCzMYfAjr52ETF0JQMBN
vJHAunpQ60LjVbVkSQzX6hhVbOQH3tOZgISkRM/jIxVYsDHQW6g3Jgv9q+mfnpTeL4jLD+zq2LnI
9tsjnY48+n7wS84zjC5svjNTMSy4c0x79NR+7qWWVFQdZDqaYYofN6/gZGP2QPDhPucT7TrvBtd/
jHNJGgOQ6ejp4TioXgxJuDojapPKdU1Jv3tv4rKCVIrvKU9sO5GNDZJ3IaxH8hEyPlw/k5kOF9RM
umMX7bu8H2+G8o33p7uRDcHttAXOc3RmiAavZTM6Id5CFxov2YICWszI2/7DOfxksGVjwLwJ2QsB
a64wa0Rksr8VYlxwF6um/1ycr/ieyD0KJcxPJFbwx3mPCOsA/2t7J40VH7xq7Q8LLngNdh/N+gjT
whHxiLzdiHLqFJRYesrueQSNBOuSoxaDmPyKlQttqTTQZYZycu5sRc/15vC/YJZ6rhh/LPJRx/gA
Ci10OeY/HwjLkaCOM3G0+w+k2CSyvSnfeC1jYNO8X9LvXYMXJGR8fEvDOm9YgM1do8CwnKWYDPiH
x2HC0K781+9RBIVdCSWZ9xMND3pN+mDXpXpxiDC2xCeT6tO2vG6Hr+9gNSV+uyLLzSruV5q51vtP
OcC3Lu95j9xHWejN8303F/58AWQ5LO6WTEV6HROKkC/10MiNo0LbR63tjdnr8neGq6ZxJaqO/YbK
Xu3zUR6mnKWBbEU3PYCUEwU0sXYdHVT8LuBIq/DpuJzh9Mq+MYgGEWn9cfwfjrNjpqkJp0whEHDY
Qn/IkchihlmDDAK4L1WipkTrDBnBks38kRtess1YGt7ddrsgRkrqdkh4q6ljnRwhKrt1IpK0FAcp
7TolL/fz0tayE248iCACG1Zue1hhOAQ2zqeEFiL3QoF9OHkFgJvef3vZ//cYDkvjF9lHLV+D4s6/
D+UaJznFt+iIGJmqFNtUKkC4F54+Et+18838qylGhsMTHyfl7zMqm+9A1dpKX47Qt3ZFytUAv9wK
dzypS7k9W03mRgu7ncNF+ATWRsDHQL3iQCybRlIXFVN1d5DdrLx4xNV0kEHGqqUx+x3ECnXU+WpB
N+dSk+/1rkfzOE2T3gf+o8S49f6m6j392XfbKf1VQXX0lxGDOWWTt2JwH2OO3/rpVpJUF7ATBSFl
J+3Ubr7guGzG6L9cp+ja5BWYPrZXttbcbzO1a0E86KQA0vNsEH/KQgv6I6eitkXuhEGzLK9ISyTe
3uZ1EPeHdyilSL9m5ohvrVuGBnRmRPZffNVK94Mc/bkE8ZXrL8BXaj9Ga9vQ1nnDcTJkSOvJFjco
h6wsI2kNXWfqUzhVixejD/GVfZLAknfPL4fJZA3omSmKUcF9I/ht6wTQYfcMtprOAqES7APJcHCW
qRE7a0VlzngSxUlcp4fUPk+qw2ma1Ft1olOVt58AZz2dt7qERTTA139O29pEsFnkhUquJzd+DhPb
1CSnwvPhpKe342aToMt5SzXg9uGEk+wnsom6q42WcyOcyuF7kaCxCY5bD+B1qmx9Acuts5jaC3DV
CDf2Lvjnu9DqPpwJhUZMW018fEUh2/FC5JfBtypLUDmWuUrJQvQYMuXUKuQGGAdWpPr9Paj5RF/V
90y7k7RFACyClduS+xgeVrMe7OQCLVuxtbAx/eWnAdTURlSdQT5PsFtfFx1dnxA9hmirDmezCZPf
OWPW+gOW9ExV/OQLBrEvW2vpk6zzwh/FcS53Eh2GeJceBOVQ4OquazyZIHA2SWggPnQuSxBryH4G
2jKB+meUHqtdxsNywZTfkzwz1yvbw5r30Oez+NHZZNmTspPsjPbTn3+XEG4rgZB7rvCPfyft2ZHZ
ZBUddeMTpHx+ozk+8EtWd8cbKgfHAl5lvdSDhcm4XERyXt/KBB/8kbqRpgFp4a64ZBW4oWRKO8NA
TzAgsr7Y702IY5LV266AKbfNfyShDJtiApIcycJsLhwD8R7PRT9IURUGOzh6AsONMk75M8b994EP
sEOg+Pr6w8TqmAJPQ8bdVWWSYwei+Xt8kAzH4Oz+TZx1ASpmV5T9Ilkv/LKpsQGMkXibpHMyhv5f
JkadyOA0w+W7OL+KJjsVwAJW7r2wvFe0lk8cOVJm/gOKwPI2V6TiLevjVUwCyQsxU4FfhxL9cuq1
li4/FE425Ks59PqXpjP0cHMJs9kSwxJKTK27pMlaqZp/nUBTLyn8PjC9HUkttA2JUKm+W2EbtqQ6
0m8J9sQmxBfhaDTWib0cxrtu759B7qAZegUXE0S01PNalV6FfZYL/nRa4rHkmpho/G7WzkLBF4WA
ti7yRRSXqxDD1dHFR0BN9D5bdcPzHAPdwBH5Q4Nnn+0D6rJpy0CvqZXqo3Gi7gLvpS7C5mMVRX5E
WQOZzDMo+NlcYkjVfkqNhEWUZJwmMETwZBtUP7oKUmXC9MvTVA8nrDQP1oXtfOow9uAxpPz74S4B
eJ3FSu9UwpLwdapd/maoNotK9oXGTDWdF5Wj0rzB7cO7fhFAebG+OGV9vgAMqGRnNRH2iqiL2hUA
8NetUY+G++ntJdd+omYRuYPQ4PyHKa8+kSyrWtF94HpaS8TvErKzRbDVO308AovCrvqZTbKzv0s/
KVcXqDTds9AH3Xqt9KVo/lCQEWwylwk8Ceq7he0ECrC1fVIF2ymmmAHj8ycNFHJnClP0VvLOW/jw
o+m2ljDuhMqsrvIukP4KLDS3CfL6mEkwET44DdB5AtjtApO2bqOer+3FAxNbGViNCHpAf5Gw1PK2
VtpdCdxdLM2d5EsVP04GSIT84ntR0NXgd9kbgRbxlR4FJdARyvtKheCb3c86gqvYwhMAyzwn32rc
iDCtAU9y/xeOScQR3+m+mORTUncvaWareLulbzFA7Ah01rtv/Azjt4uKJ8Vy1gLtMZsM+3a0gazw
2QKNemLGLXfTeqBqOeJD3dXEQTc/XL8chnptED8MmTkdSQUkLQ8HBSUa5XLSOZCIR4lnCV0Y7aY9
f8mJLIk5/+kz9nek54oC9tJ8IAqfAX/+Lwbq7ggOgNWOeyA+MYF37CL1i4aA6jkfYN17tm7MP7eJ
/SS951RAAojaKkBh6RwkwkuE/y+QcKw5YzaRyeE30wiHg+uLdTOJOyDJUOxRmxEO8DSRQVRGAp1j
i5w0Td+VTJqW8O7B+PjjSUllrzOC2zNixGOpdHbUUDjGFTyywJ8wT7c+vqRsq2SKIkKcSexTnrqQ
uVWYPplZlU2wqxInRg8OGZNrYchnglfAcTPfINj5dlMj9ybFNGp8PIvkVuzTuC1heeZfQi2eOY7P
IiZvoDBq8fEVuFy77Qo6FSeMytOmtgBK6A5+i79yAjJn3OfrbQ9sQMzyJKZvV0Vj24U33ijPAy82
2vLffvR059Nl2196BSUZEDWWOFvzTMlRqK9INmKfKbGlqCwPKPO5uOqQkf/QR5Fvf9GhqIpK0A4W
d9bLTKVhJyUoQMzkfvyKuKijPbYR/sZrcvDARgg1ddf5HHp+RytBExqVIGDdZtiDoBvVbneXZuLD
N8sONRo2nyiHcTayk/n7GED7pOHMQo+FlNqtfIvsUjzYQ6ebdLP0IKw50SzGIHE4TOGvZ/FRzu1u
48NOdk6Fj0WPVKRYrhA2NFTZ2II3F87V8K8LZ7LMhUaLpWVEUNYpfwlcOaY8ZQkaKAmqLDmb9OuJ
5HG3SG3EYmL2jltpJCDP94fikXD2JFOPYfS0nn/1skMo04d/z+MRLXLMArAj8KAOmr0DCQPcmbDt
z8fu+703omjm+xDv5usuAS5bRC4Kp3VIlwhDUIL4EGmdMvi4P1lWmxPS8ItZqRAnZaFWIt1MIhNm
JgA5BOdgLav/r9dS50ziffKmrmP84ViycvXJTE1Wd2RQ7XgB6/0JWrbaOOJlpaywlsVVHcjNLt9d
niDKZH9Unfyk1ZkmJbm78Eb2pOF8Sw99pbsNKEtdrUUw+9cfqeh78uDvffkKUYAXJ4V7/huJuyNN
FmTOiHajYAFJZCZJHpB4XgMspkeCC/Eaw/b13KT0xFTtMEozEoZ/rqhmYycx4+AqmxoVT0HaJ+dG
S1BFv+c1m9nBPSlNKoLDzh52Mc4krrW4J26+7nzx3902dZgCTDC/tg0DYv1kZtefAlTfsSVOTXj2
+88qSuGJpFibdeXQqyayh2XboQhWbAZQDLfXxNukg9ZAe1rG2P89b2zTX3GomH7XVnvmBdsDA70R
dBGlIa5wZi2NLWrGKCBS6pXm8+zNjvXzLft02HAmFHpey+M19ETyYkFy+kCB7JefNUyJiJG+TVWl
OQkf7TS6XxVyV/O5rc/YxcfKcQ7uF2PYvIERRORewqoIRP2bqpgTufF1nMHMQiROIm5mySHkAxnQ
KRTh96Zr1QiGF+TGz2DmUZwaVfDueXq4RFA3o+WBj8xU0b1lgi5j5n0rAu3wNJZSQxvN8BD9F2tP
kAhHRIL+4guurZpZxvFYvpco+TQMfvrAmVyTBpwfMWLGAHqv0n1IxCcJ66/E/nqM10biSVFQGyZB
X0cQbolb9i2ZXs74zItRuoSDX/Xjr06NZIfP8fZKHKVhns97YQ1zJb7hsLZSU3IRjk6AUJH32bJI
uQhmqYcycEtzpzi+IkhVGl9odBcDE73n8XU+GJjaRHCCF/tdDZyd33Ja0c2/sGU47RSjFRLGAjwT
QbiEptGLtqI216tn2YkuRZsYnSL/F6XgqjpFacvjLUSPHjuZEQgbZRsRovrpYDt477olon/IGehm
b1eGkiv/qpuF0XfAYoiDudRO67MZf68dxUvlKQ9jdMU5+cIaFbyF+pDvTXSpOz7EE0fBTUrb5fMN
bLyfvN7IHZSHU7MxHvu4AVceebBegluSUeqV7tg8M5+Yy85obWI8YVxnvkofNP7IdXJhCNpi0QgY
cZegghZFv2Cu4OcC5PYavecHJgB4V8omjB5WoSdw0tNyZcFcr0UhQR0CmZzRJbYxsQFXH6cB95Y+
pmWBsfl4Vq+Qd4KouxPj7YaQMmkakr2lUNDMNSSn5zrtJjmu2kWio1Ju/qjGfBF4KOzrHv211MFK
oOEQKDstYj10y8o+4bujHsoLr6B552YAZpRTV5IXFACdDh+oBfXEeCF2Z/m7hK9nyMkjrU7SvjEh
CIud36hbg1wnckT2O9Fy0sXC7s5gj3ur5N/zfBvngbeBL/FOVbJDunM2t7X+pDU73a38ruV22LuP
zVOQiHFbK8OHDeIUpGKaRDKY3MOmE+alB7rY+Wb/KNPrF2BfGlE4nfZQHuxeyAnVZwVG4zzyUo4Q
QPY5l9EhLWl1Jkor+WkVyJZ/5u9Iv9w8EFP6UcO86z4bMbzDjHn6yz44OE3VadC0d3BLeY8hUFho
EItuqhaTOP9+NDkeLIW1ZIqk6zvessm90JNi2GOKA4nKir9Adia9OQKAZX1eNsZ3Fi9pf1IKFIwU
ffOWSLDq2lZxbhXiOHo4WVxzSpp3TQZBYv9q3FVTXpp6vZsQK/7CvipNJlr+CYhneP5+A1QY1vJn
2wv+nJCb9qk8TmSk9S6EwVF72DhcTLq1bYyFIJGmsRCWoLq0WVthtt2GbODPN4fLRLQJh71IhXkj
x6Z68j4CrvcaBYMf/ohzHWjbsp4WRzSqF4RgWdVGKxv8rGq1ZmZQay1gf3i6MBjiJ7GrAJT51KhX
wLbXhQhxh64c4dOwmVgVo/7KY/KtluT3iunWYW72PQyq6X03EgohVzpJqYCBE0KL+xq5bJAICN2F
xJeJD9LcsQNKSRnMyUVy3ZkQWWDmQYitUulYJBVG/yUHy7WCv47dbDNfyL594m44bmAqHWZP57gZ
jDoG8xIvJbqAxpIeBlOV6vYpLD8mkC56KMOLTkwsM+494wIWNZIkj1tiqp/fmiNLAoyJ5WaW4Yzu
Tjvch6nnUwA9pX8A/Td6mCc6yaIFrg6OCwZ5+d1tL43xcoXlbU04mbNjJhRquemW2MhbB/fHE2tz
tshHDjEoTbngQgO9RrdIouIc/4DYcVzWJKtWMBX+zF05CvdYo1n9ZMqR6If0MBW6hGkvZsTuYaXM
aKWjd6oojZN0o3kgYbdQzvAHGyazQ7+QMTKHPbW35q5NONWAw5OokvxzwZ8JmWhbgx2C8fE6KYrN
/RMjDtwYSQ3SZviVfQN8f7RnUt6cUT2p9gw7XK5SxIDmlY80NTd/zMZp/7cRDs1Um6WUQn2WjxR5
xbHYjWMQt5BcDblrCC4GBo4KJ3/aGc/diS9m3K2ofroFgXhRUAGH2Im3Jm7qsYJnam9sdy5asrhR
EEUdSUcBN6x2nbwfF8UGDh59GdNUi5pUBXB64eowYLd4S/kt3VTwVPCV93qtO45k0CTXrA0YBUzK
dSLNhbwjpV76lFmVl9wIzLZmTHfP/zG3k+v6WNyuUo0LX9EyFYYWmtWOa2xeY0etwu5VHNreb1oP
fqKLHzL79cXU+4rWy68eaEEdo8JqrUac7jW9MWad2pRR7mkNhNgbablqKqW0xm5jOLaROUKG+vQ0
AHjO1KCwAOoJfLQ405dQoNZW7d/z4ucEFOAYlScHRd1G51MNZV+RssWWzWWmM5PzCZnJ1FF2tDlP
MIQ+jZ/hjWMEgRsuCH6wEh5yQdhbwHceGvCl1Fa1zXudz8UegNw4aPZO0u6GWYuP39pB+RWXjNA+
uNnMo7ccqJmrBf11V6vTkFTbaf1vxHEEw870Xdn4DXAc5JU4tD8RxUalWX/7spHIkVfiRktxAvGy
v2IzndkGehEDvLqwZEOKuuhaJk6lGvarUFCM7FfFQ8JOdrFye5BzQK+Kw1S/pZj416SqybMezF7b
1cIVX84C7gNgcXD9SffghQhyK8KTedZvDwixg8e0UVWu6+nqfBhGPVOi7B10i90eqy5UqP6ulAif
jw6ZfobfRfmLBoxerqrhoyBOwRordIvNcTsJPnAT2trJqgEblQgxJxAq7UEc47afQVQDQEXQQBs7
VWPDsijNS0YJSWjPSXQOmmV4gvpmYaghfqacd/b1JMQWHTdNZRhsgY3oqH704+dUIvTd73LYbcEO
cmEyiymWLFaPA92qNYAsazkMvR1keWml6Iw9Q/mM0hUx0aVqRDO3gslaqkrTxWFpADpkgLA/QccW
7wxytZD4McLFCl5xwWcvK3vrHXKNmzytAlAYw4yoj1Y4f5xlvlUHxFn3rOmBtMxJwAZfgReBK6Hi
9qPdfD7AoBxPTUaLglQfDpPs67eQyQdqrOy9yxU0T0zlaF3ROjS3e2x4zZhAtHJvRIB1fvVQiAIF
EkIxaeT2PgLQqzyDFUQbQaq4iwla8l9rQ06I3nngIbjx6pSKCbgufEfUSLOqzbDwJTpzUGDN75Gj
I0yn3VjkaldRRY0Xbpari2ZMgW6aSXDo0qLi8K/BM3gICwp1C4h52WUWsuia9AmHf5WrYnhwpEy9
re8/NIy65DRWeAxPldd1RBg2TVto6tRFxRVWKs1Siy4bO2oSlGlk7bDpch04BdHmahrJi+IbzQbe
7nUS6e+Ugb7/u8zFIHndKEyuELJJ06657qUZ9PvNcGeGrzYpOoGG/HcZVSiQMC2UIqfESsri9B5m
eb+UZvbOwJ55Pv+QAcj5Ay+WD5rq8sZpcsQVYb7xqmNWiNrXV8WYLaxv3SnRQVWBUQLH5ADDE52h
FlSyQm9A9TddRxkRisKEFma945m4+nZxmcZ5V4mL7MBlVwPDJxlGDt0pFuGLUc4PSM+2RIOYXX/9
sM55OOziCph22g6f3MSty9jceZP1hUOu1Cf7W+uVuuwiXgQzOb+4pV7v7dYrm9UqcHUznOhRQjLG
C8qGD3R2ohLrbuzDieOMo6HglY5yujsfYhIfyDYMrVsLpA/CD72++x1ds49YH0YQedaSqixKbkeN
XZtcJeT1/CrYO7V7wk2qXXNq0pGVcvk7rmCQxBC+iCJLjxT9vowfuzcMswFJX5r1I5uqrjz5UdJT
tmCEnlIq3Esy0g1AdCKUSLQOguATOkMVXHVDjIKY6VHN5aoB0BQmQ6DM8IHOQlrnDENbSWqMmcTG
wcw8LIQcdMR2xGtsZJH61jdd0wgX97BaCefmrBesJAXRY1WZS2L66xcVahQ4EEnpCQIq4al+6vRO
rBG7n44rvk+vRb5bAP+nsIUI9Hqg0lgC50jmS5P4sA1jYdPuMwgb01u+fYSPaFR+ylwWzzGxX6UE
OwY63gISFo2gvrfIgOItoDCG6R2zK0ifgwtUvRZzfqpX69D712/f3rdkELnv5MmMtjBSXZXdW99c
WaYzxwd2SpjNwXTQ3rpN3qadov1NPBk0yExBcP3wlXUHY3ZwCH7Z0rBuO1+eVlTESswQXoROQYJ9
UTlJH4CbBO5waYrIL2c3LswhhqPPjgPag62EqNhZAkQkGprtb556hvaShtX49hJJPMYUhj03pNA1
9vQ06UTykQaopr9P2+r+/UNPbPnShMn5h1hKMmW0nLjgTMwYbtVVpm9lZUUn1xsvLCpfeK3rDCS6
iz0SZdJEL3TImbueFo1c/lZPPopn5aHsOfdwL6cvZkMa+9aOXmFHjnwyQ0A9XxRiycBe0clrLjSA
AaxOA06Z4pr2XFYWTxre8gAWecrumukH17FucCW2TFNUGDZS4FnlruGURTdMs3v8H1hFrPIidNYy
9Ly9bnSAdchSKz2yem7Cssbc6NQotUdkJf5XKus8XckC1+nhDsgePeVWqH+oT9G3RcnuvYUw144C
3qS9pQ1Xua++u6bwYTk1YWoLpRz9lc1tMlQkOqUSnJaRQI3cgDcgaaxuStgHmsAO7n9S4Nfu4zw0
pfit+/jEayt98if9eh6f1aKJRIXjsZeWBtp+PQ4WL68xCIla2uX1+/Kx+NZA4d6tjg7/du5G/N1g
k83WhzIl99YZOQ7YHBmiCFd2fT2+7BE/i13nhyNlrZpnQLCWx8IpRQ8ycUq/evu5Q7aJL5/6VtlT
324TMDOhQaSl5rW/XlPkvPC4SNiE+dDpeQKI+HCfa+qylz1vbg6lyxYMgIrxDNt92Hnxr2CjOa9T
woz7SpxrceV9q1w9lFAvCip8yv3M4X4tDW7+AF3kfxQ7aMpeB0VJCq0s2cRVD2Yh3WNTT8SPlTqY
HladmsnrXMMWRcvmYLON1vA0flL/MmQMrBm0AxuL1wHTfBKzP2R2cvWa8j8yV85etWNGbfWCV5uX
5l9rERD6JIAEZH+tfZ9DRfangvTsVebHmtdR0BelxiXBdeqbKKzjNfSI30eMSZzcwijrtfmvH4Ha
PI6xXnDBx39TYAwaxCb6+Gp88u+FGpUE7OJxQ2rApzBtF8MgInUuWdP+zTZafnrlh0BijZWe+I88
BEufFkMFL1P9XLJ87DcGpvPa59wQQ6Na/WIVVyS96GmdIat5xp6YjWyDFy9wpzeAKg1xIrnna7Tt
WYlzadNQoNNPwy2WW24Q32fOo66wpNH8CWB8wM3Ui0uOQu4QA16O1sdN0sxjdKL2WPlASuoTvaRD
QiKqS8M3YLJKU2Ml0Nd/UtO6Gki8bdRHHCWNW3es9tzWbl4cxu/3zxF1k0kD3ScMJbEgLX9NhfDF
xWTvaYbtu5Neg8MJfrqmR9HQxzWdTspg4qYDxVNqL2mu8Gmecgw8NZpWqFyQBS76qYlcztJyGYLw
YT764wU/VXhW0bHYkfuTeuz+dGH4VEx+hWXl2OvCJKhJ2oLHEtmIFHPX8VimspsTwb0w/Aj+Takt
qkmpH7bhsAGdN97HWcZmgRoD0wAsH8Ajtb2H8VTmuzC5LjKVFJHr/XyIftDHh/nq/JO7aOMJztHa
0A6ECRiKXFsiBUSGw76osYTOwiNmFyH+CGtWwbDsxx+0r/FD74uHHnzgmGOwLbt8k+zI1ynXd1gi
dXNSV8jv5eZDmSpM4Tpi/2w1v5YzHHjE3PJCDmirhqeBkzXZFOuujjWAqDFk5Y7p+rlFair16ia0
VooJAZYfQDNzhxwABBrIXC/HjfmHqHP7/5/fPqV9NsK38zIyUevW4+qP8sReyaHEH1sMiACmt3os
Kn6IMkYBYSbxldHJR+ykt5vm66jsChmo4YWwzue35avsnf1rrvnf/nq6KUwBd2M1N3g5ishn8rAG
hE1KbvMh5Uk5qrBjSrUo2Vpgarr6vvQZ+4GPP3va484kLe10tqKKxapHYi615ng3QjvZud+KGpRS
/rb0aSU9dzHKu2RIM8L/kCMtcNuXzaotmlAT/w00EY2Pjg0tFFgAgkvmNbsxKsBAwKi50LI7Kg7o
T91VIcC/X9VJxNhhvgUqo/7T3CYJtzN6MhsTGkYdo4fmD4gspIPk9E9dUQupXcrmRO9iq+trx3Ax
2tXBl9inspPCfkLmc8p4Cjub78JZwY/F7FisVJsMxOr3hFLyGFcACggm2FjNlRcu0Xq1Wpg1R29r
mr1iu9PWa0R5fbWtVLtgrN/I0Q8KfDIodaB1+VicmvY8W54pehYHeOpLcspJsKUQ20wcDX0ufZDf
y4HgUcZiEBFgryF2lpBa+Mh1cPKBo4uf/d7lqLpMkWiZKQEgpWnoxbVy3F7Y2D/e0IxOOObzao3t
DJXmx8TGE2R88Fmp+UoaozdINAp+VTYm0t+hHxVilDc2bMaR/jYW18EcuMNXo3PmW0QVLV+tuMoA
Q4vqxNgdq2sv5crYEYTIy6jLrK7aIT1otmhNc3qetJHiegE6l8cCuWGnwzWcpyKql3N4zmW2Wfrp
oKcljnndyacXuP+pFpkMPQnpK60Td97JzMUq5pVPDIZOcYGs8ELjNFpDlXQGzZx6zxAatDtMnfZf
RgvYGPQH5i77e0IYmJ7JGM46vhH5Z6PpJtw+XukTVyQxJOxRvGdLF/qYqpqwMaZylUWdD4z9gzJ0
AHZTX6pcCA+BO/9UfM093YpAJi4Kn3hmdlxyEyS8zV5wquBvt0J4Y9jXUmsI9eovIz2fAEc8Lf3C
cHodSkWmwm+E59SGgftMC2VGFpP3kzAIY4b8NBFn9WiIixB+p6F+dgLd5P3eGVi9vFVhKI0ugrE+
0502HkyJhXI1o2aIeWnemvhKuC64y1WNGebikugATn9BvzOBZlf1kbBFc2a5tgfYqEvcrr1IUweO
2tY2hScKUOcY6t2NnxiFoOYxrW/cz0glLPG0RYrq/h2pDPAN8lmxUbr5R12LZCDkxKrbQcKnYUNY
SVO+BM//T7CrDgC1roSmQdvvWWe3x/QjXR3qzmvvI8GTH9j0ft1pW4ObSBwJR9eAC2lNTrXNPb4h
stVTIWA0hjysLe7kX1sk1+OLzMLct26Dpd5pJoRhP8OIIiFbaVTtD3gNy2jWzb3aMdKwr1RVjLox
OWI6wjNdO1ppBq6lwtiFGrNBpm7z5HuflDK59wYW3r7MPhYc5Xn6F0cpJXS9Vbrwcfmp78pO7Om1
xauafYoSWrhXaTPbQZKixd0svsVJZfukUFI5BbdBuV/5aWghcyuaL+XY0ZOcB9OO1fqz3iQwyzOY
DtWAEGnIvMfZVvI+WqCGkXr8kQsfEbh7rEuIx0VX+iyo/QapQWskTv6nm5+JYeLuvNAQCzw2M/33
JxBaJWyVcN8/xF2Ht34+DMPjPQ93r2wMNqtp32846FN/yoUJPOtv0upcvl5KscyQqCfGXTJjlXFc
1HubCPBvNK879fExlDyUdQpIz+nXzjZIgwADCP2zyXtP/tz2WpgjlB4+5FthKaIEBgGCPfSoHcS6
63DB+A0CRpU187KbZ57LDTI8DUmwSE8zDJloXjE/4KhBQh4WRACKFS7yrgnU9yIcapwgUlzLk24k
R55Ceww4kFAyLpC9kNAO7P/0N7BAtWJJYVTk+s14y/qgIQig2l8/sS3BsvXloW8BW+Wht0P/O2oQ
BWIpFsfkKJ/qE6pRj3gnfHbyjR7kyv+7/jfdr/cRUNZQN6P3uT4Y/cdDGxLaXMiJ72E2wo6EROUl
a0CBtS9S5BIE7aSo9a6hbQjO5fXoPPFZvm2M07h3zuf10n4lbju1hirKrMtLWoFtYAINZoenWTBP
i3PJQMWiCGFw+7zKHqUx6nClBL+Rcc7NzAPTvq80pvdB7VbDkATC2SxlmJ5bqrdYLUln6/u/mIXf
vEzg500WmQscjRWO0QLQ1pVzbU8ihfzvf9kurzfoLybBbgV2M3/eFbF9Yf9KpmItk6yGVnSqMSZ+
33T9mFs30b7Ua+EX7l96rZqcyWD+Zowj64z7lmZIrG8U4L1jOFAk1Eing4rn1n3Ioo5a2nNrmnDa
onk7cYH8jGeJu7SbdUvRNdQceM2l6SsOTKTfii9fTNdgCKV7djiN1x7+mbxGGz031cSLZBookbkU
PfvYo7d82xFko9dQ7GE8cD5n0iC/bKoqjPDHzeASuGkrYsrGkx15Uv8zk6HFDcNYEw7HAVpOFNzd
u0HPHT1TeS5pq2bZSTmwYtV5fqPGA6XRr9+jZM/LIXnBz4Ao5tOPx+nqze3B8pdeAtLbxzYpE5RP
pzLhs4HwlRGxm40HZS9KchHPcGXknV6mFf0U48w/NX/cpieorql58oCQLU+6LtkxkxrhJHVUOoS9
8e52bMvhGdmDK/AdUv3V4UCitAuGAkiEjueRr7OeFxczufFs5wZSB/JKWBj3/JNTtrFYw+2tb0yH
Ofx4ijTjhFENCoKdAPKFXwEFq63Y6Zok3QiIS+uU6c6o1bR/BeU10sMHZriGrDNHE90djE+R8OMO
n8Gflt8DpyZ+ONvMtdYYDSuJUaldm+0UcwgVFHGsh2kLMHFrV4jRx/DU8ZijTELXd/AM+xbW+8vq
viJPwF5t6s5+/uP/kSUiKv+mSJ7FGQC1gs/SczzCIawe9It7n+2BTQjJ07dkBfqXdCBsdbxopXFV
U6UmWmFCKFHKZGge+RoiTpiNH9PnTfZWraeL4j2ODCa6TLMrKCl5DpFTQHcfhpKVMnpeFnyV94H/
VdDOz2O27JJbEzIYhTw57o97OnnF8Tm9w8zq50DYtevkKpKdl7LgXI9zPzzORsH3sWK6jMWW2LhD
uwRmJeVaBGxiuhkh2LGJq2Wud9NAiBHhW9ytoG4gYzNxQToC2MpZT7O3emOHl9Yms97JQaLuLyJ2
lf6kpir2aP1W15a2wdPuji8mLzYsBp3M4ZObPZNW1ciUDTdkWbu5h+6OUP0MBY2Z0kwDai/VySFW
0wF2aqZ2uSUiRW6T/QXBbIIAMoH3GlLNxpbCYqjhzf+p35aDEhr9dldd7kdSkrxklvQ9/LMnrrWy
/KC5/NNd/yQ4E79IxjYqZ35Zc/TG1IzSC1e5MsienhSpdfKNEqVFlZOjg3RMqsgEzVmTGMpcxcA1
qwsI8He9La6Osg2A9KXby+z/Wo/qcg5/hD/8Qxtq6WbzbfooFiDkmYHu/j3BNrzT4OjZLVxp1hvy
BIamCT/OkOhJlHBR0eMzffvy0UXq7/2DCAULo/8rNzMR2tDXMOvjfoPPsRj6zsHCP0UwPR8O3p1p
tttm5NpUMhWTvUTYgBBM5/EbtxLCvp+3Z/SaUIpg9mJ8jSMB8VIuvN0tyA5goV0+WaJhxQrNcUvQ
SEYJ9imdZGge3NJ/VSlnjQKVxTA4H0+cD4fGOzYo2uBGFNJv8DX56y2bHKqwXrYm/LtIFN/QLjSz
HOW32UBzp0/3/o5w6ROaB7mC3o9C5+3X7eh8nrRvyWx5jtv7B86wiJ6S7TYlF+jcPdHAq7QAS5H1
Tga75wswmudnA0ni6MIxkgq77ftEX06B7s0/M01GwYayP+C1JDUnePJgW29ewC80Eo1B9OgzEqzl
38ZbLChg93qFGWc/Rh1wVynQUjpJ3vZnpI8leLZpWtzYg5YoVXCUAb0jSCqI+0ze+aEHlYo1G68q
SY4fK+0WBKFLsjlHNXULo4ce6njJFIGBw4iID2jHGQQSXF63j4jZWjVG2r8gAGjZEf+xZVs/jh7p
SyjM/lXkooJerpnwOMLApasw6G9MWgYuLArH7dNs1+9uLezRlQW9NZahxBJwcMDCVY9Z3Uxt5RRk
2yyzRwAR4IbsV4ZKJJaHza+PxC0HS9hy4SWzaFGSHFe+BY6K88wTm5wfLBgoQGbxpkBD+NSHx9oZ
R42qHkiXvkfvbG07+0gnSExAjN60uAps3Fsfw+KZ//cxgG79+g2IwaTkirM4aZuRmk5mydNfZ9IV
W5WPmxRNOALIqOKDmqOi4p8Xfh8R9B76/t5g4xK65xH04Z1dVoA3zgQufCeqYMFeM9Z0TMelZo1T
MUtxCilm0qeqJLUWeJTR2knWq38p+kDySdMNDl0rlCyae9HFYeXwvSrJ9+vbVNn5Wj6g7Usm93c9
rUCh6CTPYI4ud90EIvVr9HPNm9jkSLOitssc9ZhGgP7TUfaZAFdPPK8wr/jN2A0WzhxNKEAdbXaR
D9dDzgwOygR28Vkhv2t4xudoKf6at6/zqvV5cNhO1gTmjjJ21X7RPKKEJEwmioJzkmup28lHnDjh
PcZbz4MVnffgRNaHmGJJ1pciRibL9EKRw5TTbxJ3eCTjwtHDipNd3HOoCQJGMY/QuvRQg0dC/+0M
Iyvy+vpPwM37tbvE3GYiGsVXCE3VPX24lUPZ8w4FCx/X8Rkblkf3Wf5QsWsfCgJ9xGvc6JSEJvU6
i8f2qoxitqdDFT9YUygXRq5jbdITKqTvikrAIC0V8vJEPFXsFzu2aHEsw09SrW5JAsSvref5CYhO
d4Ag6bevnijas/Y8IxE8odNe0q4hm/KDHe39G+aa5EPDneyjuBToJsR87pqAiKgUnnDVPM9hKVm3
EuEyY8NGG5ZgH2OYTJuydoDI7dGb/FsTEDkbZZUiczIwy9/8YczClt6OvyyeMxMHy0ghdev+Gmvl
3trAzHNESwo/tVIVaKLICBttGaClnS+b9vfU9O3gr63PyyRMyKCPDZ3vh51fxlCHNnPFtspHPP65
ErMHSxKOJc+a3Ae3T0sOXejcPVjrao2/qkQG0ababPWINYwdWUGO2FBjCitGja4k4q/Gy6tPY8P4
/UoyP7BunW6JmP4gsM9wLyhrjxWQ5a200VTV+0xQeHWEIsiw/mdmLIm/XKjyMYG1cdXFEkd743UX
qxUUtUNoCsay6cavcbJecmfjKmdaWqyBl93LB3jUIbugM3by5TBll83j5NpJi1U1kre/nyHn+afv
hhS66JPH93CEuJO2yz+qKpN17KUaCaWFMKP9dnlQv957lCufzcvLUo2PtCNZhZlv/r7LSZI+CqiK
Axslt119mRrwtBGfbwXrcFRdneMY1KAMgiv6aKC66TxDNu/4uLgJ38X6/3HV/qPGxQNg2BeVqCMN
Ohm3s8a9HRMW5qJonOeHvNztNk0y1Kuzxee5XYovop0ExNsKtOWRpTB3leMzT6BTZ4MTvcBr3zPM
GmGLOq2mbAQeSGePBsbbd0Kkd3+kKCtNA8DRB0LETImfLYmzrYxK9+DU11OFDOGaI/f6LFSc3Doi
k5Bu1Gr2qMGjXljVGJRWbCRhXDCiMyTcA3ofoBU30+WTdCcODev6vowe59ombAqABdwpQuCCT+1t
UshT6VmTR7NYvMoPiOolnjM0y99ubaMXWFEVSHM9NVmapstd1Mduwh/SpyIesrKCM4TYKLJHrV4b
gItTEmJvRV668Jler5bwK1VBEEKTFgJRLHE3TdK5XgPMuxMwXCPzEYQYeKHN7TPMOnc5jiEd+mgb
jkkNz1+GcE/NgYDrk2Sm9x+nB+uT1pIVQtvzSZ73eY0M6XS6kPdpIVEVyg3tG1S+vOGLQdkvjYpV
+IFu/KjjwxU94QnmqaSSLUyfWaOZgHfo9+C4ZVjokgzeoi47gWqTkAquo1EYb8OuKKhJS/yH6jQL
DkzXuZohamlYvlJdK5r/RxDC7N50LvTpfjH50CQSXfuCIOpwPZuyrkCHnoPkH2j1KOUBRExm9s3p
go0xz2uVOKQakYCPh7RcO0YyvH5NVy5eDvNkJe22KNlqfBR0IcHPQ0lHQ5Rwxr8zNhiuqsg685lM
SucFlw1Qc/pG69/sc6VZS11C+swpTHXUqPgSVfAOmV7/XM30gYgVfqC0gleQbNITVmqpeVlWAnLD
4WXjeEH/eRo2S5lPWmu1wGzKn7yxkg7pV/UdB0J7aW3VVRA/XUhn4cQScPtlHGJy7PmicoztHVTX
JUuXMGL3ulEVInKDSKnevcz6u6oqVJEFGYK30OkjsWdVWIttn/3MBdjwyOQdKE6/1DXpZoshI+rm
1bxDmBlkujkaLxU4oGagDtx32uhrSM+orO/TSEzaPxQDVZaR7YohTi86fi61T33Am4OAe6/SDXBt
+MFzZ0r6pY2xEUFB0j5rjk2RV7ZAPPmZT7PxsbSmnErB1OfujJGYywOV9mryQWd9c1zsb30iNzlT
q0Tn61UXUUj7lsx2Rzl1EdPMy4K0ExtD5HyiNdfpcfDE+gSVJPTV20VHO022aff6Nl+DL89+eBsg
rpgt+iy2Ewf0XjCqGAxyr+tzHAumf/GwiMiLsDBuLvNUnZrj+PJXPEGLNkIyOMF0lsyogo2Znw7I
2+FTNjwtKL0VUme6YgC+Ov6hpGF9fiwPdfvzeZGgbtlQZpmAQ9MtVwg5R5FLbN5fVqpOIKwekkKK
nv9/sW+mJsuaNxl+ye8faB7wS3Bdu79gCLfJXQhPaIfpXK5SV+n9VkJ85bz6E7eQPMODOxc6+iLx
NNo45MGSiB2sMq/oF7/qppciehEKIvld8ZqrhxDgqMABzGl6nyVlmB+muwTsQuKRp95DD7uZ8n0y
Tj/VIh1ukIBw5CwooGQNZn6QjP6QAzGGTzffjI0c2wMJY8+dTmzBenrOTs92KkZos+46l6ehcAN8
Pny82Dz5e5Sjf9UU0hoIfdzfwbWinADUi+4S1r0ZcXdqHqKyf6craUCrgch9ncehtIVLSV0deivf
anbwG0IfCQOFBJb7Cu+NCO7zDPPSf2rErEmbaxo8Ruy55/yAvg5dQdSYqmDJNE0lsh7wuz2w2FFA
kNOqO+HYmTd3Py0A3MfBRBYcT6Xi6kcF2Njmjni+n2ogs8zuzAEOfYVQsLSa6hHY4FE5ZO5/o7YW
wYnLkYI3I/2LRCWGJqdlDMyh3LWkh2/SBw6j27d3+H+uXIPZkfesInEkLokh3yE1RDNUAFsIleXj
Thf7PQZne4Bcn+TcLR8XuTfCcafFbRrY/zmTy6n3vWr5+LikFUdAAKzuMO1s2Q5uRmx/kIMr+pVp
1JrMlbTnbyZk8fuserAeKfoHPT+KxShu2mfq3/rT73j3QWzDM7YhPOkhMkASRN+47ppvEq6R8oH8
OVHBCHGZmFX8OPS0P7YtQAkauEeqHGSpqw8lbxwRS3TZPrC/5pFqR/8M0PZxsKvnG7I4loXYk25/
bsOAStJRE6j6Xzpx8XZeC6BNWsSVMTHmpa9Emn2Yiwb29awmopaq+XJymGPELON6g4+qshYbCyzE
ekWRjKo5t2OUKVyMrD3WIAbi34SxQvMxYnjYrxYI5yRlLra2xuuAyjang0UT7zhwhI4BwLI0u5mT
OdF1UJMf8tCz6+wPAx/Ti8AKKlDoClnwXI4WJeQVIRN/g50VOnwQJ/ee588yOC/55qUu6MfJSu3B
ehK9Y8rUdgBRdNYQ7fJoEpclR04ul59Nor/WyvKft247hci5wcymrQ9oMg2A9v64o7r/LVM3riwe
FU02gg0gcwuV++a+JMcDJJ/BDxNBQfJUJSvlsByinmO18WzwloWa7USuTRDxS/Z8t2BebtRob6cm
w5jq1OcBbXAC43CeYYmwcsTCT4Ej8rXsmECufHGYLvT9pq7X18BCJpxvKX/CoAwyF1Poa+cgFz69
JEbUfQRbCfOBy9xToThKtE3u5TxDODX/DicWw91G9m+tb1Wcs4FJJrvW7aJMubuFKtQ3l8Z4AZ+T
Z762w+ucwVTi/ksFDDAFh3Dcp0BoYSnNEXaNy4yNfcbacf8eHqm6WfASba1ndPxv6oCJlXh2nYuM
Ohqhnlb/ZMfRoxkBbcNYnoheeCXHw7K7YukStNOBg+tgmk6rZHWq/Nu28ArcS2Djk354NEtElavk
1WqHEH2ys/wyMoatv3mqmEyRpz4OIR5X6uHJieiXyn/iuGavKjva/zIV0S2XBy55tmvMmxMMDDW3
x09qeMBjnT//Uig6dCtHCkfkhTZl4b3E+YBj3n7UrPmZvE03aKKwUYRuHWfCbjPZ5KY8cWL09XJH
1LF3mjf9ApmApdjYmF3OC6UAvl3wVdi8tqD6He/slIi5y9G23LLQApFpUefSl3xKNyzwytNh9Cgd
b3oBrwoWz2waHvB432J1DufsV+EgSdFNII/aZ7mTjO+NkeN3ISLGTA4XsLZq5Q2Tpx87/8emW21Y
MSEBalJq2zQ8ZHMZAcWanGuJ0wsR7BdZizdeY0ZNpdj+EKBgFGk18NhVrVd0MkJm3ciPHvuRtZFy
djv7kyNDTc1tiWdJIBzBRb/jrgI4Wems+l6cJk+Q8fROTbWpoO0PrpqJ5BzhSyP0dF8oAjEGxusZ
s4/e450sChznKe1P0QH/tSObzmm4u1IylzaTUbFtQnkXqlQCWvBPWYgTH7EFjgMi2SIbNUxFoh4l
CRgof1xfkopdUEqvmwW85vlPkpTDR0JXlw5U+gPU5tVqN3piJTSGM4ZL+lwgguAi/a35PM3w281q
VkxzFgYl2WL815hb2ywObCSw/dDb5NhrljNSpWaUvd14m2KrU4Nhg3EkCdOEImiuNJ2I7bqGee7i
p/p+PDx/E+eiTp5ssJjpEbYsstn8UGmXFcl191tH1N2bOBAGSwGFEdFOAShlYcQ5I/CbUh41MYmb
1iOhZYP2eywHuv72WP8GeqOTWr+H3gfRGR0chnzoJEkm5JAfz/Bj/RkI/jgpyLbekIwLIXOZg1Eo
R5cnIQokjy2eTVWfcgTy4r6KHG+Gm57rD7f97R5PU+PewXcfx0QmiINqrYCZikqdwD5VhHB9LxBS
ySz15LiEKmoHXF9uHIk1YON+kypdUKKhpUTr2VoIO0n/Wypeh+SgtzttDH9HBsV3SA1Gjcz8WCsK
htQyeAK+trBrE553AYxqdkvV9q2RvKGCi3bXPKNsN/2O9AB64AcQHckX3mETqyrkolfohiS3GY+W
DqWv1DBPHGDM5kXhC9i5epbTih3xakEyDoPUedifwNGcTPmo9h/bw23lZar+gzmceB6hzRx+scRm
gkO90tE1rKCSoQsaOg16W2KnSvvAKCPWIp0+7eRN2cBtkr2bJ4Wa/74AS2zFcOyQEWLmUHKwuRkA
Ua/bitnjvkROkCIOntdltpw0pQWlPmJ+dEqb4QZL5VN34wLLgwr7jhGHF8OB3U8WJuMt38AzujM4
iDXeZd9GsQQdezUvsuiMnGoorChen60VdvC9+nMDG6/VwhQoG7cXfLna9Jwcf9XvuuuNZ/Aiiyy3
wY2oZyUuX94ML8svp0JUSxDANDfxwmI6CwArF7rmbqootYHsd9vXPVDpFFdbukScpMgRZehVrIRv
AO0JAM7bQMgnkufibSHvRTYSdMt3gSqS1OIjBchm9q8YaO/fmh9VD0ZxPIT6WHuHc8/zL0IGGZas
Tc6/m1eJmn3ZIAgVM2yH2whaB67iya1Gs/MrdR/Uc68sOFYaiRAVudbfkEoXXJH65s6bkQ064wjU
qolOji/yNooWX337KNdrrubpxBEwaU5osZ45HBoKMk8g0BQ0DhCB3eZ5dqJ1u37cw/wPFVLePrev
lMjkJ+itvTKH0fChOOY8vnhZVlokbNhQnlgEiz2c2mOUFkdxB3CMi93jhiDE3+cA2SdR2RXDr5T4
98C9QHhG4qXuKRs9yFN4GGYSHZ6P7xIXPizZ+7vMlRZyp0ssJza2JYP6ZVf8WJhL7uxmB9DNnh3o
2/UPZnAHsH3h76TqPH0xLjbXupXDNCMgnTkEpoYxmxO//moJuGqRm7U0V+M+gECltcF2z+YwLRnZ
yuB1IY0IUqJby2QSQgvnpltSwNF+Utzg/zPkIb8BMz1OTvbOgsjC7/n19/FeErHP+vjnFlEZbSC5
M0zHUm+Lc23ett6zkvhG4RFYLPcDsZ+DPUHEDzK5Aj5IsY1iHu4rXa1iiSCVBB27eV3i5rN2ZH/u
jFT53WSFnnHCmDp9xInujsuXNYAWRr4V5+ibAkoSchBaDoseUZiUNJb5A/5/sm3jQL9eJFPDr6hR
zZXvUvo/ptOriXw3JUi+A98BxYyA6DcMSVHP3UyxYkLJXTnmeZn3zJjExsAuYtUrckM2NlQg5yag
cpKQutz8sSSU3rdCRV3/B+6AWObPmx3v9V0Z2M0DjD7Q3ybeBctf/2DZSwvL6NbQiCXcJQfIhFgb
NbRCCE9Xe3H7aMNwQzQFpO3XtXpARCNRCzJ0Yh4JwtfTwTtpPTS4UJ14ZDdqBElO9VTyXF+5ajLN
+duNygIxXOe4NtqFOIjolHtPCy0iNOapgYD03jDgtPclFVbc/3H14CScL3msgnSiWyrD9t231a7I
gzm/bW7iigtRu1K4sGw/2xwMK/pmQCwWCrM4TP+2nBBi2fmsnp6DPPFrRuKTih2BIWsMfHHTVwN+
U0MqIayCiPNzCsVKSwG1sddPu0raJLuuNwzt/SZ+2tpLirgaKR2N4m0iwSbdekSfVk5yRdzBrlL+
gQA03Kb9DBYDxM0xYHKoigEXSDRNk3x/SJ1V/dl5KFpiHhZT1uy/hyfJhbBd4/i2BtwqnwyPttIf
/O0lAdYE/DwhZbZLqYvaXnV/xDh/QjK+DwobxHU2z/4H6dxupKqCc1WkDwDKnAXCt86g8KIm2a3/
bytosFovkwYsJDZVgdyGKpPedgmXiPH33q3PCInx1az1ISqU8fLCGn1u7qloqIGatHO67SQ0Dyrc
3gi0BP/pm+ZsjBtj1wsv3x54zj8NyP61Op8xnDwVGFgFhXl896CoJAbiYKG/6x4zqHo325/I9zaF
hqNChYYAve2UMkB+wLxa2WvDRu1Xx0Wld7I0yp/D3iVKnd64ZEzB19K4ZYPm14dJF1j3Vs+rWD+L
4nzhI+dMx28czWf/sGgLbMU9ZlIYLAP0P6qDnbWh7ajC5DJ4YQwUbsKeprkNhLsy2oHqLN4LV+h+
7EO2kMiYfoKSGKGX37InOPGPw2y/s5S3sFnAkNe9GZcrzDxl60cTdhEOgneKZiG8JoEwg4YYdgyT
hdrIT0PRUnyzX3QsM6RxsYU34QHgESNa7wez3iCFv/j9Zb2T9zUDR5T8a7OtQa/dLDu8NGx6MYOs
uTq9XBoJGxr4b/cb05j9y6zW299B/bS5nJBBOHfrwi6ejsSlTc8kmCOD5fU07uca6aqt7PGMIac7
lQMI+DxYupUDTrfjWeEezuzC/Vg3OBAn53/0ngyDxY+KwodFStmsQOQtu9oa0KfCP3UMy2cVkZJR
1VSAh+zVousUl0bUqXsB8kGhZ/lo/hNh1ImZm7jLpkabjct1M1bNt3G5BR8IHymXzr/Lvz+GVgbZ
VVLBg2Pr49to+vYwMRmiYSxdA8/0F8fzLK5ms6uAQyPo8UFJa983nhnMw5hj8m9d7j9VmPDO/wbr
2cQn8b7scuk4a9baQ4QUcaVNfZZXUjQENWdu0SmbYB2IpMKRPftzqVKaJR6930uLznHf1ayXCz6r
MBlbFZcmruQnVV4HEyv0qlkUo/XVjj6sFGlngTyRtqkuV+/NF1/yHG5T6jhiIplPZi78F1eASTqx
lLyw/MVqsNfCNuV9cruR3B4FMttf5qzCUWvr2h1wGcnrX0iPotGlUa23nJZ7+9A7IJcehYLn4bdC
+cMoUeNtLxcPjOSd/g4EDVFwmtGugMsblnRpvhSHv/jZ5pDwSDqFDERcO4i8amomkwUdFkqwHLzv
s05163ei6Xbt7QM3/5fvO1Kg1ycEuh/rT1jU7JonaMCxmWmT5FLPYBG88LTJOnNNSLMhbQ3rGDRM
/DBqnBz/XWajyl5qlVtkjZX6KoJAVu2lhjkVmUXIAJBoIuITkWU9kFWTBl6fVDPJtbeWwJ9pWVxB
xZ6JGxv2ju8CCI4FkLdJUtQbYGsOpEkRQ0L4T2CZevi5eQ/VyBIJl3+4bpyqsu936ZcKVUsBm2WL
9HxGuGXpfzQ/dAE9zZEVMmYr1x1dsGXAJCgSBLe6WClBfNvnWO24PYa4LMH1Gdk6ot4iEckUPyIi
2omZNCPvYw2R+Ef3vPb0qJQYHGf2IMB99sRcMg5UGhY28eUoJqFOVRU+DhgvJrcl95aEwJ486ZJs
sENUybowNZ3V6GErYazU0YyVP3Fts5l/jkRSHQummWq+r5PL1aI1E5f8ExqTfahDyLkxqd983lE0
y1NLHVGSaJuULX9xWB4Tfl660byzTfW8+qM5DjOwFzR7WPKz0YLuZjyzKktNSnMrmDucikSWqaoU
EP9Cf4OE5bPjxfqKvIUtSTR8XRfjujuwAXfRiY3VypugAJGeH2RPk+ZrBuzrhOeoHcT2SGzBDhbL
nZVXy7K+oRrLqn7thmDFn1v3hUJ8flLz6sRFatNlL/4VUllYghWviHWtqFTCIlLwc+abEjkunQnY
0JA18QSoHaKO3keT0dE2Ls4xAy8rcQSRHrzixnOoV0NrYUNxxCgfw5XyZd35pN9Ms278RPi/HOJP
MQUgtD5K5BMXyQzXm2OrKeniR3ZrUE1g5+FWlOhcTwj3aGhaG03RRU7vvPRRokFO7dtvGN6dQ3wf
BIOKlLMIdlN/mrvt+7CMy6kLdAEK5JoNx3vRqZ3WZUtxxHYZoL8mzkqFHWzFptKlhvHR2paj8KeG
j1VhoJ8DHkZgTliF/5oqYGTweBLExEs0BWY4mziffTjoMPPK5iEuy+/W1V8B8bSKz9r/sc6jb0Gs
TpO9suKOzeamQIJKpRiAWhokax5pvpNE7njrmmS5UIMjMebUc4IC5oy5Up4Kmz5eBMmE0IDRQZJz
6XUKh2jBxPNA2KlbWtoIqrGNnXVK8k3L6Ln0o22phfTa2688MiblNZ5ptpUFRPq/qHqoBTyO5Bya
5W93wCP7ythpYAe01CM2uHVSekKVwP1KB2/dnnDAEI0Vn9B8yxfBU8BtFctkWz+i1JRrYdwfoJ97
X6eWVIy++G+8ZueRZb8JShD64ljm4KJfzvQDhW6ruycibOLUvwniwKCOy8bAy8L/CJ5QZUaE3Ihd
hP1GVtW69FqiARA+2SVuRMfESCFP1G+sEgPfOBtHAqKIbWwJsO2tP1nouz08tX/vbWrdYrnbdRgq
EOklYDXCaMFXnFmv/6oLq42tgyoGCGe4Stkmwnmz09cyIdx+Y6SNjiDObLRLE3hkvhaCiGmF1FyM
TrOMJmVuztwzkvJE3gCQBhlf3HjLmToq5sAakoTsQFDeBbe08IS40ZjDJ9VRpvamj8mCFl0AidBs
Vut+rlF5nfRdo1MkDVa8cxvBEuKB5db/scxZKhnOImt1e+QzpvQsyBPYRVwyswOvUZGVjjK3fm7b
fjobFBUJjd33K9uOBOwIVFqj5S2axJ4gG6DI1EVYGiJBDSDisimqiKhHGAXkps97CllYzVpJlPwn
iioswvhwi+1uur29M0aczFqtXVZC3jqXHsddcFZAWp99Ci9SzZciW6+nhhdBjEftCcjLcbImzHsi
0hjmKbTW5jWHrYbJ3pNRibKeL5+cZuD8uW+BNR6ghMaTQmrpQzq6FowddeRq6Z4ciZ5sK7cKjFLj
kaEsjnnbp8wvVl4i94mIlL+VYqjpwvrNQ/F3BcuszT7/ifOEM6SnP1zBiywC3Ay9rs1Ziaq5XfCj
dpxhgNhFaAaX5MM/1uJqLvVKWcBa0UtmyeGVfR8ACr2+/xEhbGxiqM4yAT2eCGq0Xc99xBE1mcD6
xsdfI0AF31DHzDSAh0fkuUt1ZDp3HaGnnAA8iUZek7aVDEBHZekec5LZrD1N7Hw3Vd91wk1ouHhr
x6JpGXMMu7fnlZ7Losf0ZrnlXLELuJQ41EqIJH/xwBwAsjvZbvH1YCxkUmqPvyqDNwSo0Xa5zGyY
OXxXWWiV1yVlY0fN6XY8mlyVOsP6bB5ViWGx6k4RYKblt3LLPQl3xgfUOpicusTMmEIoEdsHP8v2
Cj2Xdm1q3INuH3ubi/3MtX9rFIWmRyzjHV3Zj6jz6ZUm9ZyAvdfDPS2bpemGmnpo40FKc7rF7OHU
ajiMXqr7uQH3Z/3590M9kAYOE5M8B/SrsiOXSr3ZgKIm0LVOdJjmp0nI6F6sSNL38xVPhE3MDA2b
5xXXB+bMVomZes5cbJgxvtKUBeqb7JLTZ7CmS7YxpvRhkdVSGWLjcpN7XA7n+uiCkQ7RQrNM8KWz
j5Jv7rtEfvlPBFDDmYaO2R0yhmnu/uF+0qenzOaxKgcx0GI66GCrVOwjXwQDhm/oJ1t4OBLkXIRM
EckNebpmFWjBgmmEjKapDDirI1+3poW4/W+EYmn6RGRNGwT3FnqXNPWwjOAvJcZk/PTA1o+09OkS
QsKMugsGPDao63AnlUkSRyMcWPshQHJ+5zdS6mOIF7pfxopoCHvdjaMwxFjT3xViSsEcc2JI/4Sr
2xuJDImcmCh1jC2gZZnVkuXsGwEQ3OONFQQ3+oCl+BD+s633f5MWeFbMZJ9Mb9xsZcfxR938Qn2w
lS23ezl/vH8jKGUKMYx4wGZoEXdgMEMYBOrdQsGOo9vQWH7CA+dRUezydnwiMsTtGI9P6PtW8xCc
lgYYnuTlfnick+locZ5w72iQfTVLkXwxIaTPEIXHziTkbxqs+gCbnZM+wWkLh4CP+tjaoxidkBAP
ytC5sCSujuuh5NloDkFXbF1biyjBisk31AqsCQsYv6eDVUmU0WzC9BdKm+W8w+3yHqFGyhAzYqcM
X2xmxxV5NHof5wAkoY7jgtlFHX6dcOsc/PvqZUS/vESrWMe75P2TEyfDTe4Jw1OrGewr+EwcrVLe
bs9f02u5BlkPP0sM7frXZnCS4QM5YXo4jIbUQj9rqSIhDw4n3XD98PNIi+h67073hcxw/fKcYQfW
d6fcW8sWvyAp9wX6Nrftr8eszTrqTDN3n2R6QMrcEVH4dx8fq9ShnE1VLcAeMll0JKttPuU3Eq0G
PxPOPmViRDknD36o80fyExrdAGCN8GYkJGrMEqCbZwSmiFTApTyj5XhX3QK2ISrDdIQWG8Rc8Ppg
XCwsxQqcNSqnQAd/L+yfathmBJvfUwUfQjEzmzv25j0DSfXzyDndipuIfrIJOuJQx1farcMtnj+R
Qhyzbp+qOs3pqZdOrjp279s8jVAHZIeECrA1dfW3MdHvNs+KyXPIl5QJyoDZ1TcHC98FDjl+jDdI
wywSYQi7pyARyA66JAU7gQQ179hCfkwChUAk0stTYQpqnoMvcdCukjV2I/BFPmSdeePzW6Y/6box
HuSGpf5mp4ypCLGGdTMhBbY0RKw7Q+l+XI8ZmJ6f/M6j7mSzXRPH1cXZTs01XEb0Gwkk/GPfDZsO
w/e/X7PvalUZKGrmvaVd1sLGS6PNxWISzt6PbBYvHDGntFHjn3A6RyPUkqITYl4j70poDHTzmjQD
W+6wtz14bQE+f7TT217nUSB8hjmRotkh+DPePxWjBoQ3H8V72NiXBqymaokkcUwYO16LLmO6O6GV
Xn7rBLrQKM+OXmargQMAmOpNx3bk2wtQuZjMcDavKG5FCYLnW7rKo1+B84ucugaylBMxZvIICgcn
IEYeWdw6XSR1m3zN8+DZjrx6FugA29W7/138WjS42OSQlTFldLkD6lP9t+Q3gJodhgn7n8OYLUO2
eJluDrn+4wN0w3/nGVqXcCRBiBXR/wY5MCHS+CspIjbb1eadCQfdpvwajlWCQhhavHshM5Zh1vBp
S3BH9zCo8jRnIaN2cY/vqVvM/9JJP+c4V1h26PCXS+t4tlw7J8Z8pGZ6co+FTN9FXOw235rMjMUV
kW3v0Q/0gy11c9GO5esOQnpeYkasaQaeXMjY/t6P+G0eD/AoN07syANJVNAIuYrLsqwCjIKPJGoD
hhy6TpNsTiGkxlgKfRCuzP3vpBXb1ofrVgeoURVsi+4iPUsosqW19ZqqIBJhCwKwPljxfs0+VQYj
6C6m5kNJpJsPdQWxHA+3LLVzt6U4xhJTYDUKE6KnI1U1fM/gcE5jYe2eSnBAxZMVErdQHQDiIunM
SELR28uSubBeJwznOIm2nyL9DY9mEJqTRHc87Z1Q3JfPtM5+YFa5ubN33W7pPGUQ28kcnrtIY0KV
ISQtTuL0OjeaFNUeHAqaKjsM/tXljITWsekPYNghHlUdfS3xTBR1k4LeXy+t38PmrHyvuAoNcWJM
saCAMboy2P7N8TCq12+pG4woUmEOOw9CgzHerQQQAcLk1z3gwxddcAxfa6HTOe5P2baiRXvoCSmj
tXWnuQ2GpEkezIgyH45qsc9Pc+R3XsPFzONL2aYLLO2m9x6Mp3VPlUTBZmF2HmRg2d/qgX1mI8Km
x7YTSWDSJZtIbUkEEixvxClbD13An3clXwn5Cfb5XVvuai7QpaQ2RF4uXVrncacrxKQwGm3N8jJP
UroLjs9htGl7WIirIMXOZeiwt89bi3PxGNDPjig/3ZK3DedSHBDnwsOHwDyuun10knpS4290wkWI
CWuBrz115h4yHH7oER05kD/N7hkOcIo+UAXhbtrUm/xaeDGo0fdxP7QpYe8wAGFMOWMD0XyGbXR8
VJWqIKB7tZYfoZ2WYUkPXVb3ZInYs0Xc9HD0VCWVGGYmCFY9cgZDgSBFI9ejt2WjF577AtXUsSMs
4zQUlLN0a9Z0e/HOxZUMaeU0TQrSzzsGYLibMXMcD1y6Yod0dEPd4aUQjxPppI0XUnE7lGdf65ro
X4wXj7BqOViOCb29VxsG00GeaQOAuMaAIlKlmHeY88MIOaE3k6BMKbCHR2l0FjKzUbsCBvTvQGjr
hxuuVcKPHVjSBU0bjsgmoIOferdGbbHA88Xn+c/OF90WSYNb+PSQulwWkZho0KVR7U+m6jspwkxa
jdHvzxh/iTbT0t28y/q00NOO0jkskAOE+OOgaKm9RkXUylZGYF+ZNJcnwieeFYKs2RAcEG9LzrgS
0gAr8O3MEmy6p6x4n96JgOhxyWD92LjWVtp3XGb3NFPpOkMEOsGCWDQr/7H69Ar3toQq0Ie0znX0
c26HZZB/ty87mvNlAuVVdxRu6O68u+RP1M3aZg7xIMkLFT/WFKGO0Xd0XlAZcx5s6gbFr403DDFK
C6LQ/mV5/zwTORWg3chwjTcCmV1BuISalIV+NRYpmgObPz0gxRiNwhdIh9z8gOXDDdbY9kgxB5Zi
K3gkJ/LUcaq8gP4Dx0LwUZPAeZsVWmMR14Yb4iINOy6CC3QJ89XYnIbnEIRL9GykX7QwmBI3lM2Q
s1nhn5msbXtYwBHZaf1aiois7Ji7ai6Vl21/vrdP2uExtZWB8BST9Cvaa1cIyLVuV3PvDhoZS97g
mZdoMqQKTmP4JxQTj0+/Yrwu93OxKXXy59qkFfMY7PqDRxB6JEA9id6GCjh9YpHgBFv9GYjqjg38
dDVpVaIPfgDz8i4pg9THCW/O2BSAZ+rvWt0ywkXPcGsKpphD0jqlJrQw83JjYEftxfdIvgfCaxNw
qJGhhGxWk/7dQpydvpxZm6e7b9bii9LWCXyr5sPitpAm9rwfwMkHaS7eS9J2CYlVnwYSetZRIPn1
mxKcUNbgHiPlSN5fsvyPoWpjWjc2wUju3YflRLA5YH0+lbO5bovrSL1VM2FJns4a1wfLsBf+1rXW
iajjp3AeFTr8twycWSNyy0VPkHHuS/Ykrck1ucEd41gml/Mflvij7NuiauZKaO6blSdv3STxx+qR
OqLjBbay8j/4891EX/83X51cXPuBjRL0ZVTc9P9oxomxV5GlPOTyU43VGUJmZMyd2rRhlYq6+LnJ
h5Y7eeawRD3OT+xR9gKWFHRMZ4BeyQ9md9GQ9t2jUIm3Xxhx6YeqzwnCuh+T8/+o0qdxt2SytrL9
pNdL+eRdiIMYZfIV1a7sd44rXpejh5+mbtC+i39yxiWjnNP8tHWOE7JrlMFU+AQ5KxSHtTIfkdRN
IW8NralLZjZD6CZMLVyyvoKp2ZUpaBQvN574Rt5Wq/vvwmGg/v93O2+0lGLfp1FUxA7/35F3iLFd
FLpGRywHaUr2d8KF+PaCS4YxYtm/lie5Lm61rOFWAoEQH1V1tO2iG7nxRsCi2eI7M+9RhXDgCVl+
al2RUsEbakOK8lmCsIEAcD4oGUD/8Q8xsSpZT16g2RTmbwdXu1SorM6+jq6rpMHy+oPAsqyCBMai
2nrmU6HGQajubXfElKrUqEwKICUdqNwwSSqh6Ea4mK9YVCZpB5S8YPCqGnJijch+4+bnsq4ikzL9
3TB+a1AcKvlG1vXBnqrY+AOL/+e+zu7IZRbgVQRkGRjAMrXJQPZX6/0Ohe2g2TBQEBc+mfK52lCb
2VVSA38/xxm+vzjM1/MsNcahOZcb9kxgTFT5zgEAicHD4+2eHSzjfLsKhuXuoHeuEc58tciy0Gxz
/TyFjliCE3HGZ+uKOQgB6HWXviwzx0nDWd0ppKQDK/ntV8UuggYgdqj2ABj2+W8/FVFV3qvNT6js
cVuopFhlkGe64a8e9LVjie9BeXQxCZE0N3FrELe5OZkPqq7JKIlcNfGC91Bc/NHIet2i8USRu8lP
cy0ol/raBjXpX3sa8XkVS86cnFeDHlVul0WpyjD76bMcTiZ3BgKTKqCa6wWxtyAcUuEPhJrmGdYm
98BH8QCWeYOAt3R3iTNaOmmgwnFaKB/JprFsGlGnlK//xhTGNcYg6wA8gqnPKaV0wPfPkOlwYU9Z
J3PPBUGWSZCet/oViCtgpe/OwpCe72eQnugos0tOvfo3+NMoi+kEgPh+oKFeymtVhaR6A/xNH/wj
4Rr20K9Vo5BdmxCn2YvWlaDx2fdyMvF1y4lJtIb/R5uLMr/MYhZCcyf1zknjqVIIEB+Um8TNvId5
mvXsBf22OIgqGnA1itx8oFSGwfLDzaK5i2RNM9zN9MSoqR0I2xlqbyCN2twV6+Tq9mj5WAYrnltT
pqMHV+3qGNubLskhQle3eMHHfhB5wWc21jCKg3ID0d2cSbQXcFzXfzJkmwI0rHxlq2wnxBdLvt8N
/ZpQMAwKKr2PAabTVvlrxbiNv1KlwkqRWKxe633nIcyr6+CK+94haTo4duNNGbQiH301kSMJJmte
3oPgybZZ0sfMSodYYjPBFfleoZflSl8Z6GCLVvZrSVQMBK2obLGLnBa+CQVPfU3GEK2HMK01vfuV
s0La62WuDOMmQ35giZ/xGuDrXrL7iG30YH9sAewPscGg7IOYtU5v2Lmt/rZ5sdL0B4aDWWOGk+vn
b9MsSIZq+3zPHKoe+GcrpnJMFBwzmPci5nc5gjlRaFlhqkS1NKRq77GXElBc8728Kox6FjrZkoIV
dxjYanHvp49Bm6uExzZ53ZOpw1jQClWD+2TXRDYkUvAIglNVaow9KKByg2p70wPg/7DnyHOFFx+/
XblBXoK1l0Eei48dypP6R0reKFTlGabITHZKZw6sQhUpsnLIGiklrTeeGAioDNHd6piBGYrZTwvQ
Luxwhb/O/ZOyILFe8DGDKPpc99GzZAq6ISNA498K7TKJlxFjnW8Tt4zNu/DebvZOKXC6yJ2assB9
y6omCAk2x4Cml5MpSmc93UBD72TtKOqoAPi9VA4nu6hjwfQE8lf4KhM+q8XdzBNVekBMs6jt2NP7
3aXBHOXW1p/mLziD6akvPhZqMhbmkd6uXf46lPKM7wvgMlVtegVx712FAjtmO7YBJ0g1c+FQ/V6c
piW+FyOxS99CI9a8NHvAsdEEt/WONXbaFl/pbKRnNXmdxqzgRz3sYVXZbz9RyTbYiGp11eZTfleu
Sj6nXOozNDpB/t7+a/MzJdMBFQ7yIyUyH5pFzl54Gr/tuhiwjKH1ZlgL40Py8Mgw+7d6nhqFopH4
m0kuRl2U3R1qZ2uU4mv5UFSYkj7hZ6QVjaYUTfHQO0nyCSw7ZxwtjiCcGCwhmahakMuSmclRE18E
nkeysaPJrJvLBngwg4BsXQKmfH/UZVrU09oEuBg7v1g0Cp1eMQs23eMNQ0kjER8Hw8BhcLLLFskH
SrSpkn4MQ/+NMkm763PZXZKg7H5SzuLF/mRFaOAjA4V0AzGGb1UVKZqvdz5792EboMBP3rKc6SWG
ftbSiBGuvHOtJhzSPxDGrhBa/yBukmB1XxEgcG08Vq7Hok5YmAn/CJQUFzn0cq6gcDC6Ia8mI5cb
CnTHlGdQny5SkmQnELCtC0XF+ImgRIDelKSdmbFXy+xj/VcZmFxlZyGFWsdhVMd6oBsEiyUii/y2
qUhQ6GMMmpG3ZwF1U5DJU4ftiX7zlhx+0SViS39dbKS/ic+ab8mx84dN4265vjwitfWB1fiI8YH/
qRB3S6iDFFktmrJFPHgTib5qcbfBOLSUFMcJcfQ5kUOyiddPVSNvgG9C73rN/9KHpeHhY2SbCybJ
sj/GV5TnqHA5KNJ8nupWH+ebCl+EkLNgFOfzZlKAEorpMNksCXx6C4mhMQQdx3kDHA6oZe9NlYfo
iG9FxDLQIN2ay7O8f8YbBBCFPAvL3TdEbKudY6IXu7wE1c9aG0OAO5KeZ1qQY+Ga17n63TCLHlEQ
z7dKuyyBEuc7IXhg62xawCFoSnlieCElRNWS9LdKP7/SJK5aBvRKaloSwEMFFzHIMkpgd2ENAVlm
5OHGz/LYZMHGH1UXloIFNB6gA1XG+fEQ6qzsJe/FaTafzVk9nk8gQr0es4aYxUCE3o8Tip3U2nyv
Hzfv1JlL+YHZkpDL00zZqhlMj3SSML+gxT7U0v25kNrlENxn3tu/PZckCgNAOMC4unzgUnUVbWlh
Clq5sOJYr8QWbdbn15Sa6ecBNZ9UcFRfsynCn9EJF5p8of8cu8xB+tjXNwaSL6kySZfW2KhYwOVG
st8KmaMPHOlc/UvjrrWzxxi4uJMve03BIzGhvd8wvOpIM84CV/T9ui+XAeVF0XF8i/v6/lhqRHDo
4GyAS9buhDR9oM9xJfS1yQvQiXYkDUuyI9ndUUboG8solCbikFletbupDXLFCpo3toXRmiid1tJX
Hmx4diRwE1nhgQxX9+lyyyaZF+5v74iKf6U5OCFs6ZKB0i5vJN08XZA0PmbScfA8KuEdxorsiraA
5wTMmdq7VLqnZ+Sdli+hM5NfPJQEW3ej9bxBVzJZS1J4nHm7ye9ZNWu93qeD6yOhiz4zK7X/VIJ9
DofGVFuZvoaVZm5yegEO80PNiEBWVyRErLfpipWQPS37pD/V3Av27dUUnwx41w3LmSF+6+5a6YDi
SBUN47k7But/9KW8OO1aVDJ+6LTUdqi/ttvWd5uE5k1KROvrXtVU7vUpJK/zLhMyPWBDpere11hn
JHTqJZgGrQwYVdgr3mFrIrMOx4n5FyAWRdaK2Cvwp5eHTQ6Fg5U9L5eoKn8yDBoHmm+qFgbjHBmI
aUWah9I0XiNryAk1ETQjSbH0negvmce+gDdgLPv7oxcwqYPx9JqXrSO0TjE+50GqE4aGMn9OV0Zg
x3XayKcDOKqQeI+pHfpogvcFobOZNqlVW+22knw2fx4eeiLnjiuSUteU3g6I9Qshf+TWXCtG4Asn
OWbjyxySfSa5Tz7FTVBWEJSgiwkxUP9zk/ZKEWBh7GO/x25xE5KmQkzeE1hE/lXqyrWluKnzrLyU
1TnqKk+jZH10a3ckWjXYe4obuyGe+YlvG6wwryI+tP9NsKT9wGEu632nfdw6yHfEORsJtMXf9TES
ptO3ok7KT2lW8qtorzP/ouSj2ykuKukwaMNqX5EO0yLQQx2zTQE1mEMg2xAUAAlpDKg4HOADkzh1
dXDBd20aRrQZKuapc6MFcissAM63ZqRoZEaU3LQrpTt5WAfpWBXjDqzqrhTrF5Lb6AteRXCMSkvP
YjQOSIzE5jvt6aNaQqTHFyQaOHOweZFMoYjxe8ORirG/1ba1pycHpw/2CfKpZVFwAkwVhZniCNO2
9o1iU22tPsY6MqRVpanaUUmShO4psWGn6kbU/MoIlgo/xidZTGM+K4pKXi1DsokLwh7zdrIcEEq3
UUYbyz6FbeyGR1HPOCA7YcGyXfcYEopadI40cJ86NsIJdSUGIt3J/QkDuy9oPXddlsOLc4qDf5GA
jQx2E/tUQI/DyyqH0N0kJVTifyOJjbJE8paDot4u8W8Ke6iC4uJIpFKEqmzyfOC6YuX7ej1QY3B/
iQsugbZUljoi4mTrx2oNrAhzPAKM0vFH7ZykWeEqVyGjtwmW5pZwUNmR3sM5iRRovGLfFF1eE8Dh
O2ZPlODhGwnsF3XNg4gKD4MeobsaiGlbfMpl5R6fFeKHC7r5b8I0PkBPWQTvb27wuEGuNJ+y7rJc
oXFwGcEAmwSDredbWNLs97SLH1jNx55Y5/+R+Y5uvA2Kq2WHXc0Qr9Fsr3HeWUvypZOJA4GVGl94
UFMqXscKFuARI7hdrYc19wDOoYcjCDEDzIwsTp8TTGo7jYB8p3CKUefX93h901YGxrA3S2G5UI7M
D2xiN9E+4O/ktHd9Z62tMgPzxlY93xGyvAZimKJI0nrHz9p1se8RnlyjKh6uSqjysnZUg3J0OINz
vskLkhxjM4J7jZrbfvmABKz8P0gmsnj1/WJK6sNRE4dTHy3U3csaE+Ped8MnAuB7j+DoNDa5C6a+
1KUYC3yoRAEPBFbER2aP8YwWXqRtzbLOYF0jWAjmJkvBBNG5VncKZ2GIYJo3jYJC801SAqifRZ81
RxNOwk7pXBbElZsMpgbH9z2BdnhvY7xwwrvU20JUeMwrvfyg4muc5an24f1F+Q9Uk7WAoQbZouSk
M4XALWvDPCRWawafJc0Y/wflUKXx8qviSiTzqx4gOlWXOXR3TSy4Ppvfvgrg+0phj4EQbnZmPBzP
1weHnyCu2MatbOFkXV+WCkSyCIACtgQm96mfFFOYX1vBxM5+aTcQQZcdSru8+44qr/WsgWHB+JgR
5yycybEbl9SdnEAgifX1q6NvUYB7z8K51OhpDcoyzEP1WAoez+5//OS1MsDJoMFC+NM5wlrnDaIQ
GtyOyHATSDKuRg8z7rN8Arvm8Fnr3Q01w5IsuKd+4sjW1KKorKa2B172UDcfVh+TIuNr+HDGDjQU
3C8UhQW/rgbrlqey/1OLoIADIcVYUgb0wqm/cNQrXVWhtLh8WL3qlAdJkYVfiIZ7jLVyNB+juEi5
cs75VVEKRBkStf/oQHpNYnGfUXfbFfgnuLfw80NEUo2j60nBHHxlTvu/kJdAKmDgqPq0r6aVXsJd
2LKukp6yTpcweWH46kX96Be2LxgYxNmXktXRQk+owj4g6YbE2znFm4YKbdsCLtFzNfD6mcP/a5HS
Ba0JGsUxmKMuySTMfvsCj4+KuQ45yUKWeeFgkC9RbOK27EkPvaTMzhYLLsehJz8HU/xKdVdej7oQ
e+mnFFpQ5mw6X41z5Wp9By/R37khiRofoWE+u+oMEylnQ5miSgOAZ/3xIlTQLsIADXgWHHH8Auy1
0Mmdlj+9MeqzL7IpqHSHl6zOZcUWJyE6lcPAT/4zQzNj/m1/pDIJvE2Y8f3yclC82EtYxEROphV4
o3nzsGdIf20WD6sKGq/eAsR4AZO+18e4xX0WfpfSlK7hb4jR7nFiaMIxk1vl5Wvxe7uU4q17gsyG
lNAp4pGKW0GdgVS2w/rFiwmo5wHve4hStd4yISmGbDd6KCVI/E/xymGx9cKA6UbXE4IPdBZyQxCp
vN3gxGwPhhWmG+j98HkfRhsup+wv5JK113+j2UuDKsIhKd0+HzCjei0qHItNimRF5d/6znK2s0FU
H8pCeM8pfim0QkujBhkqqo6HQLCFQlHhLQUm4stQ7t2kgWE1OrAna0J4GO9MUcrk0czBXk1fovOz
NC/Jaj7f6kanyJAsM6zyrs4QRrg15lGaL+cf/7WjK5Clyr6Jwj+NER+3/FGxa8JnYa45y6jk2lqQ
rhdzptyKAxX9jaLkF460m48gXF8qYpgaSCci8c68IrWGG+2CioL/7ipLLEAq5luFJNuyEXPZHEHt
txkqFyDgEnmhbkjf/S5bMaBhpFPgp7TZiA22kEpfFEs8OziSsjomZlJ0rdmno8g1pukiFZEC3kTt
CKqzSf5qR2CQPmHndVtZHzWIaQT7b7OVM3W2Tr926rtVeT48eMHHO6jo9wder+XiK2F+tDtOinFz
hXkAc88Vknw/jTa2ZlYd/BfRcbtLRJL6R0omtjS2YbguKVjYOgRnE29f+pqL/VI9bjlCR9vE3BjX
4025Lc99TVzOGxAeJlbCIEOie8fgprMazDpeaIgNXpHegDbhwaOIfiYBFdN/ZLs335/s0HRH1jmG
dCGUcKMgmTEccWS5NTNqHQgWT1NBod8LxUPMg+5K1hgET5HWS+/b1xcSaJAJmbHbpOXAA6Ys5muw
kzKY4XBkpGSHvDe7ZN4G6dhbOWBa2QvXtLZntS89F3M+VODYbiUhEMO+pkfojy20rcXjb0pePA9C
uPfa534y81wKkAWZb60Uh6zh3K4Kp33tWVtN9NyzdSrSj3vG0EsJSkBmvuwT+48037zkhDaduKG5
bDbnnpJn8/ij2t97QKAfGrW9r4tZxyxKAxDNLv/oqSVYOJ912USfkMTIKRJzMBx14+BvSAhbIPDh
P3D/Xn+UPf1muct0olthqvVVd/poTrTG/SKdDEwk+mghrQKyInPBsJ49FRcvoMiv6d3PlmtN4xnm
f2Wd/fepcu6xqSIrR12O4qmahXrXQ1cbK/lkDopBUBaKuRmIayFdl/XsZEZKjgy0rBjFitFG7eQN
NlsYSCsEbQmtWXpmgl5D1Gu4tasfnL07wV5XA87xeupHxV9Jm6GJAWo3sS15I098N5o3bu7MVI0Q
VXe+rViZJm62M6rjsUH3T4qxtQZ7P4V68TnsTOLMYEf1eZy29P65pjB3pY2i7vbX7l15qxHp2G0Y
qgWG7pERptc6IzaSMbs/bM6S/yOqadjFtH60oZUcdZUVwnNzE8QBd13Pt7lUGZqKO9Yhyln8r6cw
6eO+ZsqXwI6+R9nh9mXHleVjKSPGSrHkeE51Yip1wi9DFqeVQ38K2nHCBhjTDd1audY9ZGzEQydd
t9YiKIOnhBuVLi9d2EkU6ljPHz2ZF33DN0n6NfBKyerch/KSzpDaHy4BdCjd5gk6JcWFpcPwZObO
bhOcpS21UXoJu6VmOtMz+QMtQbLORJXBgNjP+KX5B0tn8GcI+lUiRMbMB0T2hLWxYx7pbvS1sd42
2/YUly/bzJccgwlPD8c1yaialW5+p6DoMUaoXsZaYDwv0eBXRVZamUCMb9jMcAH6xu43nv/GYkna
UBmvelB0mm+sSO25alNc1GewROwJiFhW3nRQwJKo/ZUodcZeQ0Vtx3EIZUPJtTiVTUo5FrAO+/N/
YR03Gh9qe6TnUGeglfZcKnTcQzt8VH23KuBYi/eH3jv8KWlvHJt0+MHJ796L5tNFQ0feh0BmqCMN
MqF8K1f8WGlZqFRnHk3UZKruU5gjUpkNpjWcwWRCGW9eLyuoEma9AjEkpyduIdpivb+5zFWwRuiN
f5JR99hUDH9z4u7xZ1rlXQtlDphCcF7V7/CKjoonEsVTJBAl7ZWJudp9iZoZLpEGLjN+fLjt+4im
QRLotuClMh5W6DrlaUQmm0NN23d3bxV8vWGPoH6q17ext4KPu+Ms5X+aMrddS0+B83EH6NTs640H
tSuz0QSQn/DVdkdYYGUX1qWGLjooA434V6l3JfEuhxgVvDbGNDmUsQiZ5H9eRxuqC76Ipz3Q1oh2
70jLiuUBIllXOyW1WfwgHkoWec251F8Aeovs1XtRpwS7N9z+T095MVND2C0bx4JGR6ywvOXuUxxy
sp78yEFOqAbf8Uf20VcUtdLUI8915l6cxzYeIIE2JbhBCXM875ZaBX6lEbiD19hGwhZIBUSjhgyS
d1+kp+HFBxtVGM4PswOaJdfWQWKK0LGCsiTMidx7NGPFXSYMSqlX/MEZHllp+/x//WPlbfFSfhMB
CVTaahAw2K18HDrOaldfU7YhJvCHK2KVC19S7Xz19QcMDPanHtJh8cp/3uiFBXirLlNuQM7dLEh6
/EyKflkNFHOq0TKgXn/UM0yLViFngwf68hSoIaCwt+usaVUBRQJ1qC5bSfr6BIWANrl6YFbXG81b
MwiJnjUQ8I12rQ7G0tOfMas2/+InFLCsqb1pi1n7pSrvylAyrZxljUoZzCm0/xAvEEeLKmI2C9Bk
CmgObymbpnL9rBouUriYPy57nSuvDiwW3XedxCp6MNf5crPOGjQKFT3JFySiEQaHrlstKguNyW8P
dMllc2+X183fF8grelpzF8ziaiFKbD83zNRZKGA+lL5+LS9EO6DpUdxJ3HbKhpc6CZqw69Jq8K3u
ckEDpm3f27cI/KV/VGwzNIGaZZzXcdjGGTxDF/t16Bj5QjlNvwEzmiz+DSUv1HSHtWB7r3+yp63l
MyeYQJjIMVvAppTO/TIcMyX+MjteRzqKf92rC8FPGDXhQEkik0KwiLNwasFMLql4SWC6vVNex/kG
TpfelrKzMHIuJzlJ1En+RU9GVAb/QOazXtnFIq3PePuggvEE4gySeswgOBYAL2ulbEWSmzOAI+kB
JIGJG5HHat3sHgwvdKFixqtw2E8Sgu+NxwKnccn4kl6hyGRnbtRzaOrM+cYmnnqB4NGw8LKocHcW
VgmIIWqjZ+DdyzFmsQa87GUwvo24tawUVqTZL7cWBOJ9cBy1RSPCJf2YQQh44qeDaKYwsa25aS+z
k4Wck8CWICtVF19TeIaEBi9O8LtMEFroCAy71SJNs5QSBC3MYtPGXA4EXOH5Bv0KBF0H1xtTcQCR
iXyDrk5DkCOZ5Xs85bBuq9N4983u68Zoaxo/snBSVbaERYlHm1kI6EANwHeZVBf/oM5QQUwupQQ5
vFmmOjZDu/uMQ96NN7YmmIZyG9GeiBW6okdz/QRGzFXCCHMJUFgtmVYWwvW/IdOm3cX4oLDk6g6P
hkdse0gOsH2mHvGULg7KTQ3bNSx33ZJUH633Vz054Sy1iul+0neOmRW3ATfwB6maJSVd+SOvLqcc
0/2GVKnDROd6+uvWfDBkBVY5srvribi2KOBAQ3gOIjjLruebk/M4Ds9Kp0BaEg+iYV9TdLih9qoZ
g/kkLvEiDCcJs2Li9ys6rJqixo5qDYkAhMEkUxvWuAQyIl2IK5ePdlBQcTGMyn0WFXL9MIQ3qdKU
441JdQalXK+5wpKMkHv69q+L+xgR7pb4rzNSRxuCP7TzyU+iCfoSJpoQltoDY5QjidFZxCQ8Moce
9vqt4nIUEChNegvYxHuv9lo4T+Lkch0zN+d+UT/IO0l6a/Ag3lbjaKm0YTLUWBAzUtUQcCNaz7ac
ztZ8VPk8WB+H5JyLdViBT7vmcKQQIkla6tKoTH2lEZqsLs0vmi3k5xl1oyJiXdgPG9c95ab778k4
lQh0ymfDwNlb6GHVolPK5E6L9D99s0JD1JemwKRko6RDmHNZBIdt1nFBrtX7jp9yfuhKxZ+9yv9F
K1rTxP87L4jSoa4CNqz8nZo3kDCc+Uj4+UX48OGi4yjO+808uMdDiKybasN314B9vWTZHkVu7pYb
uXPJFjl+59Fwk3BG4nAbFBVXBdaY9XIzfWTdZU/POxbTfpAHXp4Oz8i5tGrCeSK0qxmE0AaMEXTn
NWyMuXcYW+OEZZ73yoFl9Ye6cq4EliH+wIFpYOoKfJmQKG90nQp2eTlnbMft4K8KeT+1CZ3vCRlg
1USRqX+C4YAGtW1fk8WI3ovMeXAupImbo1X210YUcuQA+riF4uIg2y9DpFoR1pdZ+y6HOwStUoND
GdGAguTpdfO7W7gWQOi6BDsF9dCW+0OSJd3EsPv1uNIT6C9rAlsNlCdEUtLfXodTODwxbBtTJgSn
nvljRT3jsZaryvus8E3hjaDAOGoNGfc3DO9CPuuaZs7G0kk925uNHXQiorN0Owswg52WTYU2Goyo
xwbnaHA67m2K/YcErxCeMznI0zgHbOOfg48stymJwRrav+X4twF7IgwsxU5nz2Xlp1pNBzQQ9RIs
A6aYSh85jRv+xeYvTiN2acj0gbnpbQ9pzeD9UEw063QfAElTu7SJnMO5rGOzSza+qr8CCIqJaFZO
31Q2d3aw0MXSv9XfINqYJu3YwqLA9Ah6OGxbzVef0w2VwBqGZNQSku2sTwNPxokR44DgHZ5K5ERl
0504GuTocIomCReNKDI4If8TbD0kiCUGseV5/yj3lw7XS5ipN2/ACu7MVzd0UYel9GFA//h2pKZS
4twrOZFCt1kOiogQyhlAHy/JQLp+CEKEQb85cqDR+GKIodzdIYgI/DKq1m4wxld9EhtxH5XNn1/8
pi26TpURR5jmIobkshiuA+pDW8aa5d2ScK19X2nEcXJ8ELK7wakMnyHDqYAO/TkqaIuCdtoF+ydT
CbWhUqJTRzO0laquBCLN/BfFCtiOhusH5b1LrTQzfFCJcV/a1wkPdadDssnzYEpsCptH2vknhnSK
AcbU2S4g/sw5fp2atOBReirUnhUr77lzi/LXi5Bbt0r2SOIHl3OCeVBUpLIjaHeWZv1Z8Wm+wJd9
7628GOzAqkbSxoJwj9/mFSMf6mNkPo7by5DQSUhyNLycfCok1xIkGb4o3ueOUbg1rQOkHOdPQF07
T6kw+6Hsxlvj5XSh19olhDr11hntQVSCtcMdA+NHIZLTXm1kGiC1CiEIuQIkQ6Hth7afI0RAbJOY
Z9Wv4AdZC/NR52NufuRhkx61fLCI7BgmWiOWnNBUJ0kOrCcn9LULt6PHGOLIQf6BHmzE1ry585h1
9epJxijJ9AzdqbFT/lmUcParvU/0K4m/n87+KF+hFQoca1mW9MBkvswPyXd4w7z1muMAMWCvMlwn
vNaPngaZxjasa5eguvTAO0qMWDnocn7yGiDyc7ZAmcBzo1t22NZKMuwbCX+87VniVtk2inX93ZxO
LXK8nTy/jEi8/Fm24ncTr8YLh1bqCZQ5IGugcNNzHaoQY8pJJY0/Jcy5wN81fRT6IBQWkfaPsUIe
E4fSF+Cdw+XzWcHYjk+aKUK9bU8OOl7FEyjylOGghVzKjUO/hN7UqyUVAE4bwuwC6akHqiz8fScj
FRm1+nxIAo5A+31+0KXfE6p2z0V7okLU82YzZMti/cImLBKuUU8Wdf5Sfr1FpzSBnletWD2cxDWp
IVOAl4gB51drJtvq4y0fEJZm0zuKa+i/6zmTpCPDit2fd/Pf5GxZ1PtMjg8F5Lu1TSDJEopNr8ME
zviEJa0aDooQgiZzGhshgN/RApc33dw2rxc9E7UcAlKUDsC7AJxbT6FabhxDj2eFz3v2oZ6kXTjw
pBDG+cqZAOIPpnbJtsisBz+i15Gw+xoy+McRot5FmjbynLaQnWchxKUARFGTMUlXMqg/qLeFaasp
eMIyE/zRehO3dGCQmzzKSdIeY8IIT3+P7Sd0r+XjeOf8uLWjZm7aF3KVMBZxD4lsohcVBYubMT7Q
rybW57Wpvn9Nd75ebgfs6mJ4z2cKkK5FtwtlDdSl1EJoX8Gz2e08x0gIjHqQqT1mjdxXyukPwMw5
pad8loEuD8xLHoakofayGCQ8GKZF3nIWvzz6nX1ocdvIakzHLnqDAR+idvcYUa9gcJm94YNBXyxG
0/VkOqG5u/nOB7CTxWV7M3g3EKJn4zQ9aSDWho0IRiMiVPMxaTCcoucn8Pb/qC7Ipx/19wNjH/Cn
ud3C759u1AW8x+EHDYtLnQL/LeT867HE3hLn1jYlE214ai/0FV3OQPim03KZIQZFuRR7Ybryx9Nj
VAzwbgijejSqxl1n0ax3mDTlxvdHSIG9ZiHwNt21GAPBiRA9pC13dpQfy6oR4+pJcIiynl+wAhCM
s8AmG0Q1D4e16S/j1L8TZwuE2MjuiZmUFNck1aBafmMH0ICOF8ffLOJAfabnxZ2qzIUdA79CX9ye
Tf6W5IV2RJQOt8dZyD17KbubHIcEpeFLy1h+4s5y1jZYQv5jZDqaxYtkutCeKP/wTCFLggsnscFK
JOwTy2DG15o9jZpqshbsLmzEyZZYWVEuwsUSONY6xasXcWl6pio7A0vsJ/a/Cy/VRF6Dy42ZOtEL
W4zPi1pVf5ZVuG1PJZTOu3VI7goNEGWR+iVq+7CSlqV6HWjK6C7/O5dsVoJsK92JETbnhX1Y8IHK
I0eHwJQWbyKoP7lbrqQMBzfucpaOot1Q+IDleRj5SEVgFrGXinbLW8LfsxEjM3wV9MtarEcMzbF/
8txJRIxP/3ue6CBDZ0JPsNa+y+GVLJBu4wX4HaMqsOsWN8CbUHnsYGVKYhpUn4nRtFqs2r8LPGuj
cwQe51lPB29M+Xfc2VuaFezIh3X8uc6G7Kwd6h4alDBVB6JBFEQWoxDugL0bHUhyglj/3UFAzNG+
jEXynXFGU8MoVYtfiE7cCNheYBwFzh3FrQvPQ0WbOT0wCOigs3OY2MHO3lfxT/R511sPZIzti8tx
IGi+PoMOP7iqqhAFbQ7ozizD+NIss/yr62AwWaNNd8EKmTB9phQo2MaqYFTbvWdsRvATYoJvlGZ4
hMSvAKFWdlw/8QKW+vo3tAVRJrTnOXq1EXnqWQ1HMdB978exQD4m+2xUouhK+lV/Aff6DqncVgWE
ZJlDpPJrUbugdHD1jUntOi+LV0+rBbuV/IOwb3D+HkRIxn/g70dUC96DaqJORTefdcxelzJLEX7C
toqUvRdnS+AAFNMw+fhMvv6ZQZiV2ie0ot7x8clCfb4zPjUYHdo3xphEzQ6mi9NGKuR/ugr6E+70
nsIl9eE1WbdtB9j1pJQxwBFUhlB9bt2vrIHUAuHB1gigxlwyEIPx2LIq61gyBmjX65TUwVSgIOaP
KW34uErKVSM8/cAWNKjCQEf3EYhO3ZLiZOsP7pSAGMYYvF5DDdRyTHrw24CPfdLelZjLLIx63RHJ
f5eoh7yybi3KKhBGzqmCGRb/1AM9r4pUEcv4ZKymXClZoCJtg5/BsW5UWzFVtMMaUQt8AB+yK6Lm
oDCsrjEhFmlTguj4FIHUkap9jhpUPod8V3c2gB8b3vLchacT4kvyrB2xpTIbItpQjYYCgji2Z/XD
Fbx3dDs26bad+eKBxIcl67LPQNqBxAqrDv3+NNjY7ZeJyDEMR5B9AJli9p1wrReq93kCtWAsbS94
xkVyZNlxCJfWSza4qwWHNhcly70PdcEpfepMvVOzPhj0oKcK1HuZoU8txICkE9Q2A+4Me2VGW4FT
HdpQUOcndcYk+sIBfKELz+3vg82luFaZ0nDEzUN895ovxVOV4HdCVB2ZXBniHhjV+5U81iwjajR/
/SJizeorx6h4pJ/bt9exaoy5Rc+2w/GLUkDPiGFO7C5uxiun5mpPl0ejWSUxy6G93DstukaUNOwz
r0EvRuaFy69RpqzL9FF1f4JajXosqCaKghHgwewHPTKw3qyIgYrcxrZbQ9VreLJ5pH3Q788ye9Eb
2zajbE8QuA7YsAsEIPf2mUWzVOHDmzGY9AUeKAhvNy+8qH1lJq1B2QRfp5easJuofv3lQB6MXvKP
JX0dkAds4Tva8muHhKE7l0kaXvkwuEITVGHg3empjhSjBc8jzN3e/2wjpsDn2mHkcOZvkzR51gVh
33kX77O6LfSbk5O0CsHS+7rxf24pzJoGFOFHr2B2hqp0cjsnYzjxn2pbX8lEhZr+bNWFi1qzlyWJ
sYV0QJFptz3rZc+jm2EIWUBcd4Geiw6E4GTcoBCcLj+vKrfne+vQNdP2OaDes4ZUUwPmcX8uion0
F0NO0fuJRV0S8Jcn+nwzfqus6hNT+xRIze2KpOqTfHMdrIWAoosDDOMcK5M7a7+jE0BlQEU9ga+P
HRBX08U9YfMkqTS+NnbNftexMFCEDIXpB1VWKEXRjcA1vLMS8UgIoysyUTiSOUGphnZVIAKFz3EC
PVWp1uZ5VpfuAunmmky5EC0RAowH3eObPBPBSFMkBb95FTOEDGcUn54uIyhCPpCJK5Fmgjvb8L9X
o9/Tur7FA+BuwuNfvAoPZLRQxhT8jYfuOzcz+sMob7NJrgfV5gA5DKxmdSU1nvMwr6arBIhmoqim
+843n0X+Nnm/FgnhpSSPyhpFNntRMXYSfEj+DCO6Y/TfbHrMLWlPzCIRMj9B7h+jIV46YDj7UFom
uwyA+F/NTUKsb1LWUQTDxWnocqrNRE7AW45hhwzI4j6J8mXI2fWccMm2uaAK0K77axNxhHkmtiXA
bKy8LGBBpYMgQXBwqJ2JKBInjT3obNg56IZjToqmx855xKdYdjP2j1h2+NADlc2heLnftLRNoSV9
I8+wc6fN8FzDMGXenW9xPtogfFNiToNL/atMEnIVBdul4s+7FtmMbFoc6sePk4MckjZSQYh8kNd4
JTG1P+HlnD/pfm2BS2WE7AUKMqZuWmXGcvkIJXSkFoofLPdB8wsBhE2TaPjiqO4juBBO2RbhKxxg
HfJCI6gcCvxbEaYPEU8eCLDKWH1Kg1PmMdvpgloO33lmh9gROEqJtv31Q6aSWFijWgbPvTmisGWT
doRBXsbWv2pivv9SkVYKMWHHZXa9hZBjp/ouKHTTBuotl2LtG2ijbcRevFCuQovd08Msg5rYt5X0
pwolneqHH92vHq1wHhT1KrnBCALTuaZuvupaS+dVQVoOzSG9XSNmwXrYePG8nrTHhVDX492XAcxw
M67Hdn0JI4oJ7QBs8wFI058c8zqhwgA7SSQH+iI3O3++YIoEJcSWz2/NLzMV1Pw/wdlCgTVjqcXU
dOEiQlZWybcQeWq4TblFMmtwYtdQ78WRKDZaRkX8FPWWj71sM35mN3zZ2yerwBEFe/3VJeCz2mUl
3aDp5VYIWozj67MyPLsfFyoSRuNjdhRCBFu7MJm0ByfjNXDWx2bm8YgkVjkv/SD6SfkNmG5Cp0sm
FTTbAFIIGa917UnJrB4EUOoFYDdPOhhnJmz+dI9nGuL5IHA3cPt7oTzUlv5urqezJZK0yyscWxKS
4nKO0hZ308jX6F0V1xkMDtMJLg0z4Yl+WxfwnTHX6ZDKAK1brRtT9vY3D1UTRFGqCV/tGIsJH+ds
HQ57cZcjV/MR/xQvhf8IkuXNnAqQ54dM22UPpCX0WoIgTmoVpY8AchcsQ7Ea3Nedn6Dvse5HFMRt
vdDInMx2CpcqH0a9STYoFlH48Mk0rTOjnjcgJfTqQnaDPQ4vGb8MqFN6kcpXIxDx1NHzpY8VejcN
df6BrE1XW0S26mELbDFmby6giQ7eFEF89c9biwiTNWhLAI+ghdy10LleEKfbdiLAIssIdhByK8q8
w9zb+p4WjGYaWlh3V2ygI6hL88bkOlo9Dxk60xd0f7tbWBRgRqWmuF+Au/HikpvAjBKQZpHYrpaW
TySlTdnW6Ck8uvY65C1HhCA+x9uJeiVqoFeHnu+cdiGG0SMSsuQB/5A9vf+5SAjbvntUJ7J8XOm3
985+FVr+xtDFB+fkrgTJL1BJl3Fppc4LXMGGtn6b3JveCd2CvEPWgeeNWMwVLZBv7C3M6ePUk+gI
vr65hKQF9osXvtdRJh+PaYBp/yNWlqx+ed7rik1R3wvvdDNIwJBjwqbydTigOXbjIbUiQSS54xSx
Hk8AmkPLm//3GIA8viiGOHVm4tk07EnlgR91YZLwm8ubxtNxdyyt4J+V5e2Ves//BkrAfuo8xKfG
ksOuSYNdBwQvCuvrS0aNPlfK7T94UPAaUQjrci0+Cq3ExCuQY7p2RzNihdybkCRjVrE4e5bGrGAI
8XetytzeiYheHaqs1vYGNYbeXNJN9f+pzNvG1sPAK73snUtQh8Sa6SrlH3GpYg4bZ5NN90lzlypd
AnDlzdDBuSbACmTtSwV3pSSwv3ES2m2xjzRBVwrL0I1UPfIyuX7QLRie4A2ukhgfXi23sxOwn9Xx
mUKLoBNelkLTdL1AdC3LT2l3nIMbXoSHDyPVJq5bxzMau5jSfvwL/77+r04lrL9CvsOBhTilhMUC
u4DYJMFujx9Blj4VjQZuXNGjAg+7mt+d5j4x//I/73QqHNw/waMjGeKopO0P/DrfmecWTrlHhvy2
gzhJQOn8Tk3U/A79yc/zpabou0yk1aDQWKEf2lGkjEI1ojG/VRZcoZeCaLUIGzru1t6Yv+wLl+wn
Bf887RzUQ9RqBTD95vLna4ohT9dz3PWdWvvD4v44Owv2PuyQOgqSZYs2xzbtBCnQtuOdBGIoF9wL
qPdcKXZtesjaHbYBL+ruK8zcHBShXxCgIy0SKAs6YekBuE7P1Ucg42dcNtJ50BkAbYVgUB9uW57A
7EkiNNysXx7FL4BTNPPjMphnUSwkXxwaJJtbInT9oAOBDx55zj8zbnb5Ii3fDn50upc6zckNKgrM
rUpAhmvl+i6TLL/M/AS1LSPwFeHSLqr22TYmBdsXJIlTfoGNgIoqqfFLUW6qPcVHJLn7vQ7UUQE7
qRpS+cVs/DD+g859CNKn1i5B3mzTCSaIPRMXsB/WSJbSS5X0hT936ZxJTUU2cPhEOCEtd+P6VMLf
5WRBfQHijBiTFzQgr/JdUdfW/5EdwXNVL+5dXpdR2IXiJWHLaGD5XuoAfKApwU4cXh2n/iiDWugC
fq5eIaCIzLwFmTlVd6fAWolnxeLqIviUguTodEmKkn1A8XpM1GPzV6wi/HcFjhKS4g9Lx5dN7ImY
UUQ1OG+XDyXITMuwqTQrEwRGd7g4SqfFroAdMnmN7ZipTmZV6nG6W0XNatUshnaHjqgtvJBpgV3u
LcQjiGJidbpqp/64mgMS2pq8t33ZNak3Gjn0qj7jOImnvM9YJ5zvsgYfhJkgGxnrLdFEieR7HlIF
CX7DRHyAfcK80mORBUkVRcb7JrK4vhMapWB9gqpx4OjLczUBg9TFT3ghP1bCBUElDEHLt9AHitZR
I7DXedzckgxTQVxcLjf0QcK9l+cj2FeWew7CuMpQXQJZADYg09lyRuZ1Bl5Jaa9p3xgUl68Dipwb
Dp0nVCmcb1gN40eiG99muGtuzq6D1ZqgYZIQ/YSVc8msy+3pfgJTZqnT5/AJA6VS1eES6BBWUUTR
cykBkyd/zmiklpO4KGDrKQY4eVjBwKrlkiQT1ZncM0Kqa/z58XiYVB7eUzJyF8VOZ/f4It2eULtS
90Y/N7/+ZS2xgv7ZQvVbFdR4iU7ni/Y/5Z++jjTLVYsgzfDfw/5n1uJRTJ1yi1A3jA/agdDIrTXG
DAKJeAJI/jDEzvOyPNCv6wH4FBpO/JdXAsex+CkVKoUYJxbdybYiH5+QGO3NpBKJxLTVs/G27Mwu
bHQ9oGxF4dLpnaGl81gXmSxMbsYWwDYLV3Wz1h/zjAoP/gXi8RV0Xy/9UP7DGgSHIWQXAq2AEjp+
tn8FU5ZWDQ/JEr5bNQlO7X1mUxt1Sz8dTvIRpnGw+1SzopqmC3DDGXVE/b92vPgPSoq9vTLFeqgU
/ox8CAJiGTVGkr8lcY2wRRnWtaqcw+NV1Zc2fWCle67eLlO0lgxnWPI9mxJQ888NV/Axk+x6aLRl
/YVBogyuENgebJLbJk6Qel5NR7P2thLpcKLQK3PNjyb3lpxn98lwZ1NmOl81RUYD94viBMz0e51C
IGPWpSqDtSOUObEXVzV2hZjBIW0Pz4z8t1YeyvYz4PrI2xop8ThMgDGSSzUWQFthlG7dvX0t276G
P8GAjf4UzshG7VmI9qExsic72d6XN3izete7MYoIFlXlZ5Z+Lrvk50Y6otH/lfvY+s4uiXBhu+Ni
E0tyTU6ElgW1htiuPVYAj46U68PO371L4Lcr6akO8T8KqwcVBpUNHOQrn8qt7UmjtVlTBmRYZIqM
xBj4uBG88GoX+VcRZ5X6zbfCoyBEy5wkjtaNkiOtaWWg8ElbZkUKYnhpj5Qf6OMV8TSAzY0kh/hp
Wqx2KZheSpN2OjhG2C9pjHU3Q5Rls1ZGr+o6RNW9BFH8PZU25rF+zY3zItDqwZJ4ac+cKsHLXjwe
jyCtvRbnTRfacf9atBSH4z7/izxJgzSXomFRe7ljlxTZp78o0UF1cb4yMZts94KBViVW7SkX6rbP
gjGcbzK6H6pd9tybOoaKlsTr20uvpO6l3jAreYLGDTDPgsnJZQT6RrIjF73SZwqyXlRA60FRv72k
EFLYbSVHn3GdinMA9RM3riKJzl3b0iUeDeMJvwO9/RLN41lAv5BUdDaecHCvao/jn/XY1w7uOFK4
f1KcVnM9uViL10K3cw9Jowwv9mmxrsWLGZhDGg9Nwhx0//C+eL1lXSmpsczQgpJAxUN2mdFHhra9
5n4UacZ4++dqdgj8h1z+Yr0Y2IzpKYBVX1eW+MQEYWYwXPc2KQGXfHCxMAZ1eUz3hfJq2KvMAHxy
W6+Y5xKS27xQH5L/5WvmGl1P03+IQ5/gCdePlALcy4z4BlAAiNtl+EctDjE4B4AVxHWp/dUdeYXQ
bReQ/57FvMtZ4OOU/0mcMRLoJ31U8/TOFnwcvxS7fHonVOVXE9EPKrJtYBvyzDTE2IxcxyegvFLA
lqV9RPLyUD5ve2dqfToDj1wb4Pd+rvm4tZf+tESdZil0dM195LEFuPHl9phOcnHXak49z/rjhQHB
sHrLENVDfGJB8JqKSAgcY8by4HgZ96CDRKNvzRC9WA5DmEb/r42yKp6aXvDr/IZrKBdq0R6GTpHf
x5pzXQKLG+Tp+js9ln/AZmsliThl5hL6S6NWkSkoh/c3PucV3oDubWmSEJUJ/2z/ue4x3A/DENeS
n6Z3MkFN5gSRaZ14LtlNl1Fw7jnwAzZp02lhHa6VSDDfa08VoXkTh3TLZHf0TnT/W4HGiH1eqSQ1
HgncEojiKwK6roEGFVttWJRAohgOt2PjXJVeo9KK/oASqzIWFe4RgKBWFcxBXMRFrJtpS4eUbWg7
Bn78nxKQZbb2VZp120UhLC95/0k2vnlg+XMAD0iuBPX1wYpstmpk02BicxHA6uItJ5b9P44kG7S4
HixkFGBdhtXsXQTfx2upPdZ3lQGsf4AlPuN82PREbrt/NAJ88AdcFxuu3IenHfBk6UwoqgIHYJcu
AZ/5OkTB4EeimzbtGrPW+JC9HlLE6n/MChwV1tHY6Js0Jmnsiseo6r9AsyQW7QoE3KeY+O6Zkq7w
EbWh9oRhe7oM+vytSejMChIj9BHrdAWvLcyrZsM6/wCbosUXoY1YOmLkR+/bcuqTInu0A0pM6bfJ
TMi5iEO0guzuCVZr9IFYO8VbPANWzkSE1Xe5CttMgtCCS3kMbudZXQl9SjIeYT7TTWPs+mY7wR0i
l5dleAxA9hyN8o8RfzX1ctu/Uf2xQ7cTXoMVgsTqOXVDZV8hVMsAgGLDSqgkTmwNMY7so6nyGM+8
Cmm7/JADq8TOrGm0r/8JVq54yfz6STNsKAy2ZpOThSATTv2bqtWgZ0pkt+BPi2us0u4Q+4YXi71+
zAx4xJn/3UuBjValh8hlYTGcMnCfkGIRUi9z1WTLxRM6NkD5sHfNnoktFOuL4RhILXxPvFWZGr9C
/zYq1sK1fyiXe3w17D1ZncrPQbWHPm7uGTwyzHwn+y4nu9pSAMeCrbx/z0wXagGaZxEkil3jBPyq
PQA0uwFymB+y0SQv9KiF3BkghTWi5PIk4LtHc7SY1/JiD14NirrwgOJ4eZSsa8ct1uyZMKoVjQyI
b3phUqv5WyLmMpDlP+i4RPY4JXPmpkQUVCvyPq8wwuE2k1UgQW2Zw67qmAJLb0CcN8EkeKxciDDG
4ug7rKtA80M0lYmh1JYNCtuAH+DG/VdB6VSFYoTu8OT7ptzSXYT1n40CAGc0a4v+lza5xFmTe4Qa
5t2pkW0F3Kliu7e5SqtkdweubKv7F6LZU7nLY9S7vpaxOQXetDgSp6EElWayK7UgAH8EJ/rOGk8T
gIPKSLc2ZrF7uhbhklWU7e89WJA+J3ZIqC/6L6MFTd6Mjqtn+uMmEsgdLTKI6XNYvnwuCaxz4tOY
A+TxESVmZsXZPTlAg7mOQlmITl8U7Gkx3nBP+pZss3GhWEkOfr0iCqjVmKtEBv+UNDBPHfMfyEtf
JEU+A86OeOaiFhnMwnpaXn1qAQ5kb+UBRa8RWI0xkwgQDxj8MCQhHb7I/8ww422Exg6hDu6zAQqY
xNsZVKLt4EmyxHcCwCuTl3eNjiztsXDu5FTJBJJGftllu8l1Bfe2pO+65cofxG+pfk/MZxPFGc9N
1kcGghVIoBNqz9nUvE4sFD81zciZyjMc/MHKpTYHW8umNAZ2//936uvK7XFLkZOUmLPkEq3yeAqr
ECz2nR3rowV2nsbxDqLUyPVm5wilWnYzPOk0KWQoZ9Xul/QXYCqbDvx/OLd5Aqx+0JQUHlffAAzI
Q+C+HVqub350Vu0yw/rCFxo9zuTHRytCTsg66soPL5s+s28/MShoidlGl+HEmb3qabosWa/SVe2i
HKXVbvqXN88CCa++uOVqLhX3HZFfdNkj8GFwuOwK9e9yEyIM9SdH4oq9tfbrR5QrvEb9qblNHUvI
agOJF4stPmJBe+niDmSzxQ6TdEUp6mqiL8TYDlkw144qN+YFVIA0DGpc3+CyXGrxylyjYCWIkiDz
W8Jd6lJMe5lhDtPSXonHdYMv9wvY+1fnLCk/YhJvnF4+t4N/rcPBuJNCDbJ+LJCmhXOsRut4sMX9
aFkKlVV8xvWHr1K8RIh85W+pX1408P20RhmfoDZLTnUxOVHot0PDrtk7YtuI2yaIrgAiai+Iazze
Tekpqi1b38fQWtF40w8w4zK9R+JEExOs5RfwxAPFwnuIBrOg9u1NhLVpTwd0Ur49eW6yTGpSlLbI
YjW6RxhnctwHXjc1+ey/7j10hxUIf2yFD8MFUWv9Vs1eocOWC30NlC0RAN1sIfS09sTWhC7UkwzO
yGhEt0462AnpULW3Wyf/tgTKn2G415DbJJR12RDJecfdXJPfzXPjXFiOnyp85B1z9ph4XSZsGmyH
muc2cGU8LYc2RzO/EutGcUFUFB8b0mv0ModH/zsk2efWuKEGqKgAEQo7MXzVYuIkdv6yXnPpYLwh
CxkXSXpB5qvmSS83iNJVctyHuuu9hPgoWbeS43ucLXC+0QiEOGGPvvWAD8tb/e3ddJILJm38LluI
pFKCzZYa7n45PgaYptgrDrymVDs6273MrKw6mw4mBRyGeXGCYftuLf1XYxt6wY+3mHnVbhALDooq
ylYdl9KBvG2DmENmPG23NwQDY2rggJeF9w6CUfaPzyvYJ7fUO/S7+kKt4zAvIkKv6AKKw+OYXN+q
3/BGEgbFCzzbyiQGOSoKIN35bN+AzJVDchM1DHVU5NRPsGikf16BT+k4eJP758qKHe+1SZMdPws/
3DbdbjlkPzJXWddoQ8ETu+HaDUPyYVUFntLyzxeDsB9BvwIayeJ8Z00OMp2H94nfuryyn+ULGSs+
QsPx4Dqt9AzEwhc8cbpbB4ZK/i9Kab2LecB2cq3YxqDfZrALoA0ZQwL4ADbZ9KEWJUJVul+lwPYl
QX8ucfrdjP0w+DH3QSl7CT1Hf63Q//sqKqIo1J1zl0xRcl45lqFFs91TwsSnZ6dk+gSUQQztDHh7
hK16SC02//DJSHcJXjzxu6RkDxomoGGeJ9CT5fqh/Ixhz/7Ol60PdbBgZAk92DLV1NcbYJSPH5Xl
E5q5PdS912mTTcSDySCoppxXstA07rXWy53ljNMswxKhWmnJGW9ST88s8oQKSSZZHdJ1haE/oafq
M/wEh+Je2+kOwibyRqGZNo7wwtJDmmGrH3Wssr+b2fdiZ8VP3le9NsVt7aUsrcB0XPzDvcQE865U
b/elvb4YQTNxEUJ+AOg7u/EZd8XGqtZV4eNMfCU0uqwzePduCO+msY6WCuWfiwubnXtpu6SihIfn
LuCmsQvKnbJ+HCD31tFpkPHyaq2lVG+WPHBdEebTa8HNv3BOIlqhSJJ+zp6lZbRkm4Ql4iKwMoH1
pJr8jEneaFq/M7cW1CBFmkDJUShKEpJkotpOdDkRg5g45WKQLXlGbCsbmf/yjiZ5PvjoteYxwjym
mJxZFxj4cMwdSqN7ow1ybZZHV0l7Gxuz8BrEdjYH0es28BNx83dIGPJ+/517gPFvPZzViFB1B+Tr
QoY/14MSbBATug2LcBsBc7irY/xjfnH3uf8RaH+Y9RiXA54uLOoUK0cEHUHzlB/X97Dl5reGbh70
0oWK34QjSXmTke2usQxubdGPu/HOX1IBNSdUFlI8XyxnII0rC6Z6rqcpZK3OhYmnoTU09xYxbwY+
LtyobL7ZFcGDVSYC5bVRszSfIJ8jxDP+zY4dGI6XMB76KK5VHpqFpLTXormziR5vmc2QXT67ukew
X9XUY9wjoCnWGbJvmrZr88pk1ucpfHUb9Zh7ecJdJ04d08i8nYUDSLGRR7TbfUfYramELRHiLJLM
2nhfxArrDHbzXOrJvtb9NVrtXf41qyGRNrnya8EVKaIEDZS7aJ7UaM8bK4mOaTLJH/4c1AXk2DxJ
65PEmBY6KhD71A2VJgOcFMHXMTNaLfGCrwAqECF62jSPatKV1QKpP0WrbMCAkAvnlTm95TxNpmd7
FICvB9flP6V/gJUQSQ2+5QRlkwGtD8P8OBw4c62u7aZcz9ZfPFrKfh0noVGBvc8ljhaeBa4uV+2Z
ImZqnTIqrWjt0wjoXuy5jAhlNKPfX22+m+e125bQl794J5wAV3lmjYSWJ/iovaLAbVR/FAfqyxA7
KQ7ZRawap6w3QJXEf907J1Fh6wrZILo6VW27m090O+v5TVDvWl4EldJ7pklddKBCjYdCtEtqVl0a
LGGqWvYgdNkQjf2Qc5DHU4V6zpaqwhRqeOpRVCk0v+EOslIdjW2pYSy+TRuoRNAYvmrV2V95aKmb
1o2DPTj9XtD+5ZEFJ7AaT4oUebIRTwa770r8xOzDmZEYzMPzb4KQxRknJvnHDD67F2mW130REIpL
q7BYBgfYlCkP2+BOYR5YDT2ZUGspdQJIKOWXbidIRBPHM7EURuUHmL3iut5zqfvx1pWWYt91jwac
8hUWjj/Mv9TnM8cFRxGxu6cDlLAKuzYwbZYWynP2kWukN9E4OMYk3hb6UpJzYW0SRdtN1WtHaGCB
gz0tCRQYyS0ri/MWmN4NzDE42c49DFiAJ03sDe+iVPkSoYF+tj9hVnEcvOPMJIKEL/eDDBisckuz
4NI6rZuZbgRHIzJXNc5Blo6tUNHajRZz05fVMiHoa/1RX+bHco6GuSIJOM+/u5CZJIxc2homcFGA
kChx4+CNZe0Xh2W8RsqxytmNNIDwxYWGRYClY6KUtSL/lKimURZqZj/ALmH3dq0DW7IF5lZpJkuV
s46shJnQl5a7r3rU7lGb4p6c8s8BzlTP9uxKR9gcW6vzm4bUdjgamPoL95Lzi3LDXHDfmqEWU/pg
pV58yCvNBOasYCoEIsCqQjhvtfwiY8nWUBM1ZzqwIHKBzPpTcu2W85vNj9aK0FEGKUA8P0U334Jp
JIBQQ3BTdTvmY/JIvz0mJflryg9faPiNxm2HlL3IVN0Z8TdvaY3466FKeUkXXmgi79srYRW+qHCT
BYTP47oD6M0L3umQ2iFmWwew/PPHHBbyWIL2FphphAkoXaLBZO2B9IWe00PW2VzmZE8VFHhpAQh5
VsOP7uKSMw81bwBkxiMr8h9LPQuVg2/GFwhdGi9n5AyFyc7fjCeBfRdC3K83phlhbiHG89/m5dr0
z4uCbONnUTrG9pwCcsH8NLXiPWFntDUG5twfgEUaj1qK1yMafJQF+d1u1fTsaisD/PAB+xOcDA1s
iUub9Wap9jgHYbzNGCtMHkgeYbYoiT65ghSqCsTOnP/sE35NOJOr1b6eS9gVOIHXRSljScPuzYmO
Q/RO36aIsP/NPL2A5StqmViP22dUHJiOkYIvrJu0DmnMwUyEri5fJo1UPsiGFxhD6Sr3jevR1uDO
v4C4esJkK0uL71GsavCO4cRdq/mPPC3UWrBYtTVejSm7L3NjW3hzXEReLPo/dRcwsf03bmlgwyEK
xGLYlzFvdcZ89JAcgsj+HOcAyNXUw/b3SosoFv1C9iE6XxVv5rjqeWF2oaZHu+ou+168v9cZIR2w
5hvKaM8WHkYDo+mgjYWdDg6Y7jZa3Q1YGMJxGT4rE4ppa98fo5AREnEVfpT5V4SguBobd7hrogJC
Pza2lZZ0MunaawmTZQjsJym/Or+M3zSaKmObYa2JQTd0nhdOHQ/qQ1mwHr78xxqhoCSm1/kmj9WZ
W05rpZf1Fy7izkKabCl31tESd8Sije4DjvVmuw3tg2LQNvbmtdBrYygq9YUENhkdMTUdBkyvztHP
M18ZFH8Cr+Ot0QBdyirrETeoJVYTYQG39rLsYvLXGAWh8/bBB4QG6X+82fK9UyVYWrNpqfQiy3Zx
WxY3cGaCN5RLU1LvSHYw+GJJPR+kZ4wbdReaBRF6q219xm1T4nFFOwRSUZ/17h2S6xKOSqWZ9cs7
EgrU5a+WkfD1OgvPUNeX+ynzyqTTzp/8EmJd/HrPZOOoRH8oB4dmrURVDMRdOfm7D6WMdIHC4Xb6
CzTKrAgFlBdheMllZe40wkq2Uk+iuQoRk9AHDSoEl5pMY/zEKMgRG46qAZ9WPfkbgHP0LUd/Tu0m
dRoeDssjm0yAB+tnlVJSEKhZUOROcIGiDExp/ns4PUDX2TAeUjjz1AXVcEBudi+pIXfWzchRHTJp
G9ChEzyopvrMcyMAgbtEj2d65VLTdKhWDbwSlgb8C3F1AxuSxAsVWmMXLUnoKmZSxqah9FjXvnvT
FjfmK5q4ylmnmFyQNnnUQrY+myHMIo8UApRluD9nQPrSABzDcLjxaPtxCB6o0+LMz5xTket5flZM
XHKgb/FdIfYMYfyXyBgWYD3J/Dl3/CKwk4i67/D3OiP4uC5vIAAwo3D5DGTWRpCwVqllb+zshARD
Fi1m/+yZHEu/9raRk9TJAA8QJFccPpz6P8HSKkQpR0NZN6/igj4dB7naQJwmpCV8WP+VgqRye9no
CBzRSAjO871Vevw8HXq3UbgNbOhyYGvdz0buTcw8EnFDeAWej1D5JgF4VK6HoA9BXWUKqeceBcyQ
4GH+Ery+q7DYujzyQUDqOiyFdrxtTswCM9NvpbHVbh+O21F9vJJ45DvYiCbfep7SQY2mSylwSIbS
qqwZ7rpU3h5Ysvy59Ma1SKv0++WuArUqJwjrVyoEbtSZlNlSZz7M6yUmQU8NAWi9/F4oDU7/SSTB
96vFZcqykhFtokXS5boXp30KMHJJ2+H6jbYHbl3v5vH4iHwvYlNeqdMOENA5AP5S+Ic5LhzEIgIU
ZrHTMnSTJ7+u0nL55dEffFg45C4EhaKn5Y8HqbfpDn+4ialNXQBKzI8MRI2t2/+l/2nejR2FFqWk
YgR8lwDMf8wyd8qvyBtI0I0o6yFkqfU8bB76S6pBCsKWQQGLxQjrqap6Zd1tA/Mlo4/7qvZXdZm+
CUfuqTcwY52N0xfnRUeciOTJhZsQKDOinNHzpLmRa4Ar6hAJ76TkKpJTTBFrfRay6PIn4rsW2Klw
DBI3C4sC4tVAD1tI6u6uWkJZP1POpB8ekyFaKnWw2jSvX79GKiQwf7zQieFslppst9zDSW1dX6O/
Cb8+x37QkrwgGeQuInekCe55rAxrocJcjqgosiDpvdcsMPg4yeMnRk7QgCL8eI8Ua8hbt5gdVt22
IkFwwDLbFMyavNaKzbQnNSyT974lsydredLOhPhTCToBlg9H01M/GXeGEbHzPnFysWkAaXsxFV0Y
upSvLqgiAFn0RMhrm37MYVQSWgB/eKPRJR5oAPeBt/tr/sS7+0f3Fyb6N/XPPSVqrpGnfZQCDh9T
7BdY4+N8wPL7lO+ZRjQ1UNOsxzdIfymbKORINE0cjmmqX66DcZmrBBqU9lO2spQiMXooD0UUWBwB
EA96alGlFZM1HlS0KbMdYPOOpWcYXutuyugtgh6nh2CPnxCDkeQl1Xy2Ge35MFyBlllWFHvRlNCZ
t/Oenap8H1l1ZOPWVOqvDl3JKQpIKeG2MRfSNE40iwVJcTqtZ80Fs2jhPzNGYcsbh5rcrqHA2GPi
5T1rFaaqo29Tvwo8ti9CWce1N1W9yDfQA+EXkybEYVRRwa0+n85dkZMWdjLCWCUHkU9JialJsjRb
J/+WrbvmcaMmH6MXCnpvfzDo1aRX8sNN7q0AG0FqNctycy07K/EO5XhAi8hqhni6I0xWpba7gt72
4Ra1mdLGmVhZDuOCzi6a52iEf7PXfg2zkyAxicZJn4DAGFZCnYjXbenwipRdN+s9nssHsK83BX+0
i05qaIyIWThOnrjmFaUKRNzD42tUV2F02G+4bPhJb/+ha8I4bCMzqHqBEffNv3fxtYuDtNXfpLZR
0zMhUtHdzIgc/Fi43Et5xpU6G2ss6nWapm9/X6d+UCAegk+gZrarylp1jXzPdR8fqkvwnHKCyHgD
G7rbt0WeJhD1IiTQZQjdr0YxR7uvD4su1jIakZPhTv9JXybh5k5qj8HYruZcym3SZ4nD6sOU4Hw3
AOtO6rZXo3JMext0CsjkB7wtjyfKetvscq/wPm2q+wxNEUO9viCDRpeRLWCVhSAvvPablqUiG0aA
dvI8QAqlDd8YJoVCOcl4ECQ2noQwvC3Q5VrWyTjDXIe5aKi7d9lAEKzU4Yh3iERZSZdGTmDiWNv/
cbB9e7gqz9LXUZTcwZzhdbjS3YMfcXzPcWSI302g62+pT1mWwqY6YcfaIAH+cZ7c+H1EC/WyQ5Tn
7kZLCVBNnDaK+dTzbeAdwijnIIHrlGounrXLAici8xzoGLynNc117MMNVxx5RXsupKjeXwYefaU7
6pfmdhea692SmEcAVESwyANp7hrsW12M9yhl078g40DR4Q03QLBbcGMyYX0eSIzowAuymRMornNM
Rn/4n0z9lI1sTDo63F4voUI2O11lYbgwrTbDWDREHPVwroI5C0QksNSWMpYh0oyaLj7DKh8x6vm3
JegXOH++FstfGBqwnkO0GiCjO87zbPHD591ipNZ5jmk9amHY4Z48TUPhEk1nrc0m2U4BkeIPtDOD
7z/oy9ABTbAKRVxKFNOkTnLeIhPgCL90/YLCf2RQSkIz2hGwOHIGRDsPXf2bmwcApptgXz+6jsP1
mVPkUs63LyvsP7liH2YqdIgHaNZlP26ayek49bgkpr4AtKHNm5qvK4DYA64FAqISHzZs2xiTyDe4
WjMf0V835oxujlZLE7Jm1rX/S+9Jv7GgorR3dMSlhQM7gl8hAQ9cWqIZGzFJ8r/sgQNHwzSHqGSZ
QbHZ3NxdFmWi5nNuKq3z8X1JPFLJ2pZuvejJIMf8QgrZbN/hY9/XIfu1v74Vu5ESPP7VH8tb3zFF
8/XZxBHkUF9kJQRsJfaQEfAXHR3cPxcVkCUD+iT+6PV7G9zeGe8qJrgTZrEODnIswT+7LkSUn77W
po/ZTS4qvzBd2UxO2EqoMrER6NiM3Lr8eWmG5Cs3N6kse3tPpzWN7qQ8EoXXofhK7zSkpD0pbpZW
1T89YO6KfI+LkvZpn78smD5eBsrZZ7UYO8N5gjRX9AtsWR9VqtmnKPXqk1/PpKuMVDEgQFYQ6uZo
QaDBfmos0WWTIZzZEkrx8ZvJkE0in2iWY/HFXZ6LeXkaLBi/QE7RJ52iXi9Dhw51//mhsQowtpAs
qOqeJTTlZWEJ8GriZGERKJnJEla+e+MACqOilR+M41lZeidajTtqsa8zTAf0jXvbUtWyM3CkrvdC
w60E1DJa5KE3FbN54EeCYqCITBeyeF9sElk7NhTuywXeSLyqFdDfDYBQ4XL8le0ZGtlF7NO2jeT6
lzaD2C0bouURXFR1/YuMXyIQG8Lrv3Ax2XQ4xIMlG8FU1xa5ZKjmvw+ANggGM0byBV7U7rxcewpH
DlnTrk/EQ4oDXI9FP8WDwzCcqYj57aySewKTEPHQxe1CvxNV9WiE/fvU+ETX1CeI5xapoYL8u6GP
zAyYh4at8Q/eoc3GWBHGhDiTCcQ4a04M0NT/hsy7s8kFVX8ECXzGEM9e+nMQKxpnu/DdgmlhHMyL
LPOb1T0VU9+o2m6T2z+Gn7mVHhABsl9QLmqmd31WtEHb1Pa63E1RGfHmce6I04NKp8r/Wk5DsESa
+UVdOT8gCISg1dmgsup7kAgg9tzhn6+BOUe1mwgjzbj5knVfB4wSn0dOiCUsUWzBinM+ZViStvPI
TaRfM2lQZGeJQOoNEPzjkmnpRVWcmt3XS9m9fA0R2l29zDlG478zZU1zd0A/cE2P2fLWxKY3M67G
I4flb5uYdyh4DbqJ/Wff/Vz1GiTLqbk8U0PeSxEZHCaaaQSJ8UfTmQzY2iIBH5wATS7rkk2x0AXT
2je7/6UOzLsCO7a8pMnEa89bcNuF7Pla4aPY44qj6N08W/fRyvZepU9JOKutS2KKyfirfTrt+gX+
RINcWOwHXxd23wkhxBGh8tGjnQWHAWvVPZoZipnQQ7nAPm4Kp69alZVGZpT2bsz27Y9uOBA4d6h0
FERVcNtpUBjx+3wAnKbUnqlS1ikt/wUOSlipsK3IuY+LZeJ+KRx/WCoJx1Y7NRXNpZYc6FHpigFu
cLyrkb8TV9aiUnHpP2FnAYN3YWAJiUzaAJO4iJ1dGSf3DN0X9wSOCA2oCesHYAoySm05MRyL3JpG
PEW/NsB3dVYEL+C77fss1dL7VdPwkIlP1rxQH5Zu1iYhxGONrRtPI/ovEZDvB6aLiCWWEaMBgRwb
wHzg9iby9D+FTFnB5HWyOKGzSr62oUF6v6qR4jd+K3fAbFKtiiGfkgjcQjg/+QHYBgJTDZFYef/G
6uw5jUHn5cD50bf2SsdOpX9RYaCF9Gt/NPQdDQmosaR9ICak0LJntycrR/70GhzP2j3d3HwD0z30
pplsQHJFdiOYImcBAqhQk/zXAAAmxzLZ2UU+1fcI/zqoMGuuqWj6IiQ+b1AMR+IOGPKZbGeLyQFx
XRiM9e2/eL9tTL1bQyBAgNm7CJFu6YsUYPbPY8XGuN+1Ru8Bvfz/AEflSolmMJjXzBobyakcEZz1
+M4Ibz4lVqmWkYEYO8hwnNJ+z57nXgPrxjKMn63ZAR0WMbAHfArw03eGNuXRtvWg2asU6Cmmr1LO
9X+stt7h/FgKE5jMUBIuaw6Toi9w8CDDpwQYOj+8FJ6AMHQ9ji9PJ5Q5GtAwugCeT9jQghLF7OaK
0exyL33/xflkLV85IbwSdTvjP6dWKkFqdxGR00M7AcE4NYI11xNQEnJROZQ2ThxeUhWZMecEte0k
PIpTbfK2COgLEzNJ4YYAck3NBdhdjiajVJo674ModAKwJM54D+8QBhUHRi+6+qlXb4efTZVsVQcq
3dFO+qg3LzcGyA6CME1/uoojlRSNY2VcSSQFUSpuWzbIBZ7k1to4OO6jx04PqvHisCqHTKDd/u5V
j+F99Sd4TGB/W2QCeOblcv/Jb6SlQU1Gb2Zx2ugENPUVpuLvhvYUpuU6IVDJvpDx0RhHQm3Z0CJx
bpQ6m6qKxip3m0BIDYUtucJhS1JJJySeJdC3YuI1lkDtWOnOkfE6rpuz1f4fjH9AVd6WAb/0DdSs
n8u8c8sE+ijM6gawtovaKvTSZI/RMamNpIf1Vseb6b7TPa28SLBmXyHql16sRWprW5d/jtgK8oOW
vP5i3YEMhTbG8EQgZdgKEouyWYZjN0c8u7tuy8YMxNWzQUs9L8mufc8H2OFLL9N2DotcnC2qNgyE
F35pFditVFjpv54p5CpUa0GFITPKVyYuB4XAYxpde3b+sNn7B+SBSXDpvI030d3IecvocLgCXCFk
dbBALUyeVemMUhucNPJMR+GClmMuVtYI0wkZuesYEc9EWNCZR9wu9jcQ7MtwWzVfUyZva0YsXX40
kMIx9jaPNKN0InFiSBBu7PYNeRUX/xmMMWV0SVn/mQ/OmLWqWcI2NoTHSUVB9S5UXae5BHRnaxau
lVJUOhoOCiKRcbbyUeTj/oZIVjcwalw4pmXQuMNrBkNeGMzLxTGy40PMWAKcyfie5uleBObsqfiu
sQVrfly7AQexUAi3+DrsTLiEwC+D038da9qcmv4QkKCxG12kmf7BZc3VXDK3cQ2lJmdkuFCRsb9h
+mO0b5YpJVfmgD3aObJt6SFAx8NmMTlwyI94wb9O5vFuYIkKL538vw1uk1R4BDJaaL/r1FSMPVvh
3jUCMrRmTHNCBPYGWJ/rkzgwxLyM3KN8qI/LhjD0oENXV4xz+Gk6m61wCeob3bxNLamUphNGudN6
YxwWodLXDc3rEmeHGsm5lr3qR/iF9Bg6EbLGGRqwglai3c63cDJifHqwNLl57BBiHpYx52wkoBuY
gd4mBThI7gyTFpmWeir4OAuM9YUg9lJyzdoqgyQ+d12WjuzmB75M0CLQ/M/Edqp0LIrv7T/w71NP
f5w6MSjOQciFSfcZ6E5TP1WvdA8qH78vnLWBkBvSLq4QCP/u+EEUXeRnoFGh4k4NXC+Zp4CstuJx
kJcrI6ak0Eef6+ZciMrN/I/HfT0f73eBxwQGc4006x33PajUAAngeRUPPDjG9+nS4XIyjM12U8pV
mU/E19Py+o07Op9NWL8VV9wR2Eh5Ytblvku3eTo9jPyyTcCFRQSafcxrx+3ZP+n06mqY1IonamAw
/bVfo2TlNEyj3apL9x47NK6VVUcntQrJFk8pDlAvegkIl93p7odu+3VJjvCt4V0zWlpXMRu55JCy
87zTs1MK04FaLqZehqhCwX5XEAiJY+dYf82rdC00m1ysgOR9N+muq/qJ6AP17ixdx02zRzTb7AlS
0qNP6QB6zLb992/jDFHfIHfKTJ1h5U+jcV7rXFit84qIhR0CslxshHtzc1gUr9Po4KjXFI0HS7CP
PIeQ/XX1hSiCWDUv/CnaMFDjMwMb6/nEuvSCSohG183hZEqzfvoV+hgVlgThHJlxd4xK+7WDMETo
Rw4BS5LSt7SBAXZcCg38Thna3Df0ThO6bE4C0oWmOjkdJn82EcAYeNBM4Rmxh+/8cnm2MTeg5Xzj
f5nLS6BDVmAuTVbfSnfUWa0KDL9dmtdlTOBveMJwXrMhKEFbmhCCV1t1e8UqEAtRUs9LEtHbRhYP
CxX5aK+4Mii6V48mJIX/T59AmPY+GRDvJZ8clsDzfLFPj4RaLnFS1PaornuwtH/uXcINtJZS5hpB
5i+Moj4KnPksUOiOhXIOFbCJJteCnamoc5+0jnMyrtzP8n0G/wlpTQsJ4mYDKgMlewVtpfZRAJ42
b2oOiXK83SHTWUNcD3YQB1cK2KjJFvIv1jfRRD79GPhUQ1K5Dm9NeGavPv7dw28fqv3Rx8OVo6nk
814QrmeKt91kNXChv3cj6BY6Ck2eXVvV7XIxq2HEJGyGoMl1/fR8Ixoghkf5EULosIMHhGmQSVbT
mOUiKnCx1FVyVyXHGBVzdfKC09p1AnCsei46KLjtjxjb98KSI10r61wbjFo0SX7JX7yYkcmUpphn
D+VF/rYyDTwZPwqYrPcjdFIu3HUJ69iWhj/vH0s/hZBLV3b++WWgsLD3HdtyZg0lITm0nP3LQFHT
SPM/XEaIJFPemAONq5vMHWYvRPH39GktBF6/iQND8Q1hf+YF9lqxyYyN/l3OfqoKq1FAKuhMSUWj
4cxnZxTbnbdcrtmuWYUczcP8DF3MPM+mZ08OZkCsBLlFwjda+BZK4a7+5uCZGsclDhfbhI1Xo8DM
lXcJo1xId9rthD70ObDVjqQvDX1UvxWaGZBylRhXqO68d/IWeumTTygJuF9H4grBZvE9oH610VUI
XM1cCHt9L7KIi37+pFCpb58bbSj2NmFLFzzDlEUkVxeZrge/7cojp9pq9xntG5ESor7N3fahlDvX
oAShz4aSynYDP0ADW9o+bB89/Qb4ZLNSU8iABDQD1KSMQesCflx85McJ1S1ycwtiywBQ/QWOUsC5
Pqu22ZaTQgU2KPiE+6qNrVj13NdO1zF8UKNN51y5Sd+naNFIDM5OordRdOJqihTzl23dp1bKoLBf
Yk+oU7y4PmcSvPqYjyAvTGgq3ZqEoGNRlPK/xX5d4gWCuJtFQh7ibfPaoGN8Uzs+Ig8jmV41jtWv
2e9CJVXobr25/jXqgoV3khN6ruY2xwa30l2U/1nk1xgVYmZ6xITjUQNsdyvqquZ64JkeIKR/cE07
uI+d4I66+rmpGXXySDWU7EK3CVGhxk7DkRNPC4d9sf335GhzF4qcrKw3fioiznPJ5DvaVBJvQZdQ
hDSmb0z0Fa5ZwLfo1nartufFgF6nMLmd8XCSlvIXozzafILzA6Ef10rLI+1jloF1dhHGh669BzGP
YHaV69PdZR3Fn+VSQWkpK2oXGeAsCu42+fBVV8PGplwcBwiqSEpxT8Af3HwZcCVuSdkZVynI0Ops
2uywCUbgNT0cWlL4wP5M7guMg6XjIpIOHBvAx7wY2wKhrzj6IIyVE+tlEjpuIB9fgFAoyM1l/fu9
V7joe+3jBHqaPz67rL2ZC6pkfzfdRkKMVQ2k+cIgtVx+XgKv8StBTiecVdeaeos6EhIIvtumd6l4
GMgPbjH9Xg/QHtHPKwgZviZVBVhuZv4J5Sf0ql9Mc4mf0sZJJtGrrCJnXDM2aCSOYFti/URmve1e
+YjzcKHsfP68ZAMsKSehAmPlIsyhsExMcUe5f3Xh9Eaut2XxI1ckgb/lfZUpMyfcdnyKFc8rBjfT
/Hf+cyJvu2g2EEZ2R/RB0CKHtinAVCLEWfZtjvWNr/qDoxK4bFilg+cnYdzY5+6mGdNq4dPyPrhq
zGRojXOpJaw1DWMkroD+uuYFL+OtdhCFNyc6E1xJRx4+aghb0JVYRuA+FipL8+aocMrzln83MbjG
rD2u9TwiVj8+5uL+HqEtTU4hZvYrfvlGakpBPcQIZ4OeX5O1DUiFLLS/dM2mmEtwjYVoLC3ejNau
7WhICrzMqv2Qrkib4TTDCnG5DWk7JlgNa76NSFefFvJViPwWVMoAS7gSaGeqCe+YxPJGlPC+p4HK
EkmY2EEuXAl2//umnDKyJOWCSDmzczm0VB8A18RtGElQW83H30gz6y7APkaU/GcXAtoXouu4a7md
kHkfr1KBKAqD32RtlmBGOfEXOPlpnj/8fIfHBd1nqgngFkjMXfDCnAYZYA7M4hWuw2UfMDowYqKV
kH2Er2CSBgLoaqxUVA49GQpXwlKqrkXPLEm+EG59QDqsi+WCD1w7Ea2pd/Y6I4Uy+RameCvqp80A
xGWCsd9xSbkivmdxLn5aC7i0cUCTFEmCPlJtRTP8/1m2+mO4Sm1OWeTihXcf/VbP4X++cSPMdm83
ADpf9LEE1LZRKqEyssMP6b/drJdh2pn2QSbk5pMQu88s7DtHKstpMJCWKtj1GdGK2GmU0zKeZqP1
qEyk21B1mFZzPx6Pc5buE3FZvKhNLQY96Y0pgo5Z7kxbjNs+JUIozUQWWsYBTQtbdjA9Jl+K1Wq5
MVdA5afPQHSxUzZGJLtMof7kPvgxKNjpglaBGi4uHnJnMFdH9pP20jRwyKl33aeLtn3tiQuEgfZX
kk8LE4T8fIsnbUOFbX0RuO72rdiDKWBU/Yk3AGxgUKNqmmqcOAjDXjL+anjjPsrpgr4Vd+CSrSuO
nh2P+a5YCFm4dp+HFDxhE1/U/T5QV+4pTvbPjOPah0E+3kWy6ErFYDdZRSRdPSkz9X5tU4FiwXu3
XO+X0UdGgOkiYcRBO7QDy7cdGv0xlmbctNC8xdE3MPp8qeaBhS4MZbIqMlujDWLlmobNt2DU9ExU
dxjaDQPkCGSM3+uuUg92uNQtkbjO9Pd936ezUJ9gd41pRkVd7km6LGYf19cf8VpjiBSxDc4ouj5G
BEdyXZYGPOM7rt6BF64NrDNAJAw9OxNsPSb7k0wjhUqf+Ym6LFVuHkwWh8lfJiJb+qZkslr7pMAn
C5vtU/4vkMy9F49Hcx6tvoU/6X8UPkAuXt25NOQUgx2IXnHzjJV3wHnJa9YDzG+d6yiTD9tT1nSg
I6RoJLqptQ9h9oTvQMelgUKOzBxflmPJNh95CBFrmGo5NYLTsCt7QfO7A23bBVuP+Z0iJB2Kjr6y
Gg7gtINtdruQLRZYql8I6i3//jZ/idVcULodFxdk6GA+L2j2NEH+gy4v7VAN60/AsspMLn8AVUO3
oNfVgHVUjRYgqQNEAS7U4c2B7k+rG99DB4J9n34tqgMeXRmMc/ommxgdPQzhk1RO+E5RhzLN2DNC
cC+ijlOymZbmGZOKvcBrvT99aAAhm2e+DDvq+iAgUehuKqYTq8gYjZ78ANVVOEDClLPv28zz4L0f
vyge90JCr6fpvZQicsQa6u99bBRO9htVsVX4qrwRf7RV2vvNqNycD0xTph+1rzi3T8H0Au1UWfXe
D7IovFkK0GcS98lKhWizjHgpVNWr7tT2Hn034BfO8ntIeQPQKabMWyCvGJWkSUqlf/zHn5foi/TS
wYJXMyJ8Tfae7ozcCkb8J42qZeftJQlTX3GVSHs1+3UaEl86EjT/MLqKRNihjipfmhHbvaPBvDbI
0fD1TlFXE0xuVJYiZicehOSyBsp68UQnXyvLNlC4WSLhXzQakCXRZ1pKamL0I9BXlcKTkNf3/ldS
opZoKnP0+OcNwneKIY95uhjfRdZ285gOWF4jNlJM/jw/y5fK+pvBjZYCD5MqPrt8P3yWZu+K7ZcI
avfUNYiLwOm6B4WJ2K5A0hD4KZ8nAAA3vuprXwvUJpe7leRNo+OHZeR1v+ybWI6OphWCP+3yh7bP
ibJwUjDXDMeCrYLlmnC/stKvc/DxO7GtLDmGxtiSiubPlmrz8AcV1ya/+Hw1vALsEXFJB5Mn9xX1
WDDe0KG6bO5ctPfOETmF9tfVKWJvbWQlfxRrqc+h8AAFX6Rggu3/dfQuJHnla66h/ZiI0tkQiCeH
53g16USc67nUcfvOpNZZwKFPy5hWWdffdDi7Im5wTWnHMgPWZSIgIpZioSaHwdg1Lm2Ysb8JJs0u
xJ8mb8rFDtQyefZwbOsx09wC8rFV0dFY6yL6xE4Z9HThlLdnfdditQFPp7UVyZNFrWco00y7XTNH
OZfOTmeJG7L20ROU0sThxcSWy6fCQjifcvwmV804Oh14wYO+quSR5d1Kg6c4xBqLDjUSSXmzaI5v
3nVJXzw0k7lzSHrsoRCJJ03hXW/gA1zsevrS7uFlcoXB33Oj3pgI+48czK3Ws6IU1TVbih1fgaRz
XLv3ZT/KxwM/tcnao3cRxMaIVDs3VizVeSOkZkxWewfkcG6QSpduDf0E3GkTChwFVBUBkGC3OsJ3
xKZ8B4HaFEDlOFbDwUyoVR+kE9U0GX9qwkBa9PHUswQlLdsIF4dhn79qUD6ge5a9QZGxM3fl+VOg
Yfn08nSb+0ioivaBLx8Iebiyp1KBoiFxNAbvxO+lDf99fvldP/cJDd9kS0FP7bNjKgUwTYvvP7N+
lESxOeEQqqqvSnBt+O26IAsXlwRGdANrhf7NUO65l5IWqYBhTbi0iJHjCyqYBGAqTn3hPHblrDHk
tmxfA/+M5Mo81Fy04G1DS+kr8LYJbR3Y6T6bPwEot9jNAlQ1fadpCNN5IWLsU9xeMeGsvXm8Qzar
MH+xGvJU+r5YpFfJKztnkiiEqwZVR++2PTi0917mGXpTvik7d+7FV2Eg/2AkNrU+Supy2oQxYf0y
sxn0Pn+5Hzb+xd0Z08Y9y86ij4e8FYUnMJ7G9AiNrMXUO96dbhbeF5+6OWkvxZTYtRk+3il1wu4O
XBJVOmLTIjv2ahWQyd3eI8vI3IHaZ9c8cGu3nsG/Ngi5KiwVUMKhoRsViDhMF7Y0AbHoLeKO2Um4
4FsGDfgCFVqekrRB4zz7i6yC+rr5OyGlJHc7XbLRRjPdtsOg4gzxL439yLYlovhGRdSRTYDKHJ4O
8mVHqhgF9SkmV5/FGqptt0cOQJm+Rp557OyJsFllYfuELOnbq6BrS0T2piLRE4d8LpACvPmlUO7m
O1xKN/onAN445cN/sHHpGng86eptESwONX00gndRys7c3y3D4fDFVs2g5nruJvt2fxdekmTtfjaH
PgcfOC4owqdB0D1rHF7GO6NLZe+bTAhpweyTJg/z3yCHk0rOxvFvH4lzmdUCgkWZXgNWxmoTs4t/
CQq0wkvwou/wonjn9vnLndMmMSY6jlaQ0+x2ksb/gbYWkWuhXjdvdv29uZBm1Xitt15E6L04Toiz
1btVzrVFJX6s/5qlN4uPdjPCGI25LSUPCfWw9bQorPsRvgVZtnig3n9JgEiHJgxWsI6ZAv5QzXgN
t6JGkW8KDezo86wptZYELY9RGlEp9mVJvg1ncw9DqeY9o2RqyTSOVUfQz52mhnh+ZUkGo6EaO7Ol
YQFyCyDIQuiGHnnEN6P4WErhzgUyBrEW9Nap+6LEwiWhAaHMDphbClKilS4nNtE/62vn6rat7E/8
3Vxdr4N6GBAT1wO87hLiACs9JM7vCzManMJ+IVBxh961cRbD4qwj8+X8I17MA+tYMcNn1xC2kRsW
y3xcoIF7z1w9fs3DWUopvCslKdUDqIVdEGhFVqXGHdVi5cJM28/GSqp6JLNpNsulFGQPeeaeHNOe
ervDu/drnFbuVBA1ug1ckhs5FLjs1AErPVpRuFRIcaQoCdm+tror0vz7a6kEWaQcJ3A1/p9OEE/H
6665gnlNl5cPF+kZ8AJHHx2aR153MjVjppeU5BBnhlCTLplXhr+5ON8L9E7+ibv9DTHAXaBt55C9
dePhCGL/JYq47DI+u1Kgj+YMqLgOdyQ2NYpVM8YymbL+yxULJhIGjLvjK0PGl11YTRHQbAYTKXAt
qR2LzNdZkdSDYSsGM7ptt8/p7yjITKlHTK4DxrBWJL2pNifVan/OrofhRvxzYYgFKWk8liombsRf
hXCJbS+N75pm6MLJclOUQt7q9uT/JbjlIND/50W6j8h0GO7AD0LBs4SOaqjWZKqDOdk0NCPmKyd5
+trl66+HgoHz0crzSWrJVjIarudppTfvMcW+MI1MhmOQ3p+x/pbNGz/CE8qRXg2hhe98BntmtN4+
Nan8rYBwG2GD3vrrSero+f3f+rJZ1xfchZsXv41x/KYJpBFw0og4s+uImhZJrhJ2Uh1IgDh82FdK
ZmB5OERTmQ8PpWMKCNLymSl1EjsnlBto04usssWPXPYTDBIYtmqdCYyuA7ZJ7cb7hw9BbUxkwOlD
lkr/rh7lMSSbd2VKEBnJ76yqpZK/of1U79njOAGQeN0Uy4ulJQEuHvQgxPb/SXJfQMjVBr3Z16OW
00tpLEe8p6+awnwO87lyu0f7NtM2egnSqPDWZ7ZHyZzSixYJdZdrJoEby/Dz4qrTiiBsPMkPY2is
nxe5AppN1T3YYtCLXoW6K12j0ZK98XVpuBH6epF5ONCMVTTTgycqh4THekGMtJfP5eto1v6JwqOw
/VkIjITV9SJ5AGW0jjDk2eJFuIxwTRCl5g3aHIdohHrOhyeXlWFLxc0TfOjVvJwL+iU/s4W2QU3L
mXr9R4TfW2oNxRII86hn3XHLnl/e8ZcgAcpO+9I+6rwzn3RnHBdAcdYhfyeuZlXqwpHzgL+8JtfU
UPD728irk0u0613K5ojZx3QE1MOwBdrKbYGfXjgMMxGWUxsziF8fJ6lKNubfpOeorkDA2yTIg952
Z9spQ+5+IOQK6dRPVwNyivmFTzBlrrrQJvMRcTaDVunSttZHnMSaLG7t08ujzsLBt4YrSuVRvBl8
siZt8Z3XpdTD6Gc3sEE5X0SLv6BSlqmrKI1dxG2chLqjnZeGfaxDGPVmJdMdKsdZHn0zzsD3fZG2
KTEoHG3QAGWRrqXDpWyU5bx8UdKnlnWlmu3NeZBmWweNhyd3uixZu5NZexQYHcXXiOJbIzKL/bJM
4mVz7XO99pyeK2maHympKlMJQ1R+woRH/ybcZ+anJ8FUd2va9R0XeRilWTO4YHMYISc1qFohqu0i
5sfJu9QforfFsp/QHCuBcSg/ZW1XBzMUqp4Xd+JaYC7p7vF/ZeZk+aUUipNu/rbzx1Dnw8Kvy4fR
UW+NR5HkwOHjKE8db7+NZr7P6TBlgPHcCAvXG6aAshtC4hZV4prQcToJWLey8qjD+8uXu1ymm4lI
d1t3AePgl+yR2+7wGO05qi3f/MBAGR4CXKa/B/32LFOQ9UpwjYtuSCmHJvXaGLhnA3Ve30PfsBWx
YFdWpne9EOrjKi5KQRxPfIR8MukY9E+mbKmhJJVn2n3CmhVyj/+bnvcLCuoWQZkz1Bxf95gnJ5AR
3I8hmj9RVAnJGbrAgauQYs5UCEIeDjUha8GOjibqqAnWLAgn7SQWrsoQDfIlaCMnFnbgMwLKHZAW
hIu0gy5joPVWAQ+o1kCiqaEPal4uM71eIk5iKF+2tvIfWIqEweHdB+zfQ7SbMI9y+F6p74hudimJ
HybVpdpimY7Ah5q7+s4hKMjaoqBUeXnOJ0b0XOiPMHIv3uxxdvg05UgQ3HB4LfjGrHstZzTSayoC
hevTNw7yMdGqj2GRa0Z982Bfi4ptFkisM44GXPO23cf/A/eh7aeGK9fSw1/QN2ORX52KX3o/62et
pPIiXt0VeCiT0qvqK/JWiwyid1j5oijeRgXzzTiCd8RX6eIZv6FTAEUq5SrjuSgRMrFSD5Lcdb21
u9ObMI2VOSXDyuOwZe/LhCZ1lM0ogrVEcFoMIw7esegigkmKMEQ9gEGyBc4vxApOS6pO0AD/MAXs
LMozESQsFtnNJkC7+hXJk31RAHLk/RZeINbARFKUmBENw2stwuncBse7oK+SbHClSiF63hguy6R5
QeOIsVsU+13xdwsRR0uG6YxA3V8upmjddvyc3RIhzY0kyvFoGmw5H1/VNV9ncfMaUmU4W+E1MEB4
2BQHuW8xOcQxc2Pt0AoF/2B3/vvJMhEPP2scO8LcnX0F/1+gnBOWC5Z5zcCh48ZpS1xOezzX1XbI
O7jk3Ou+02+gu5lUFZ5bhI6wtv3CvToGy+75lq1QpkWZ/0OsEyaNEZDyonM6tPyh/Sz3ziqHlf5l
NzE1gQLWGEIcDBDg2HCKAeHCINbA/R4DLOMPlCWmjzM8V+2U7xhQck4i92T/VzO7sCciUXP0e251
WxLm/gQ+bFmROXNbwwh+k4yyoaoJJ+wZggXKSs8A1hyMCeVWgtRlhm3H6U4rSqpnvw2W36C2bmhE
UYs4/NwTEtw92cMVfP42M7xXCtasuP9CoO6qNWl7PBb4tgSBfjveoM9NrXmJmsTbEUYwnyFbCPr4
iu+j4d7Yr7VqRy/GsCg4F3SPRkvQqX7oebX23Uy9+ljBAAM796uJF08Gj4G4nysVWLFU22fChn2A
ujVSFBwwtxwJ7eYSrV+IoDt3Nm1vo/vuzlBA2PmKrlINPC8xELCIXY0a4q/8yV7oHDRh/GVY4SVh
9S+fhPMpv+HbpfV6lV4koPG+nFYfot/lcF0vuhs4Vyc7r3qmtVYVmPqFJe297xDjLWeAdXgZ108K
w3b9fiJvKTVTB24s/ButZGMEl4tVqOZ8GM5C8Foymj/z8bPngKb/bmAeTXmXhgOEKZ4MMINaOX6e
nQ9IeB3dEpisvUGFEijZymbd9du6h8zOE3dcTW7cjSGYCUQ9UlMWVJjm4PC6bRf0h48GWxODdPB+
XEFxxavRhigqY8st54yEv004+XAsZgJ9eQRnR+nM8m+jZUigRoVGgtC3q7aPgsOaod9k8E644l4g
YZgrBXPFPJo8Mjmc20694JJeuh72Al/sNg94+KGXnqgWmrMrH2zLTYt+k0NMpn2EtzMuFB7hSGVo
2VTtZbAf94bf2+JNqDMcRWX2zV34hwpc/VcgobroH0TdhU93nmgvuVwCWcbKUlIyfJodScxoiczj
D+7UtKCsN0nsvQsLfHFT4bX6+biy8egSgpnD4VRsI4PYOpFjDg1yjYCYDkdHo4L8WXWeeEIwGo6t
5Kf7sLBfLyq2fqWcHYpDimS4vYjNCX4gdjS5iEw6aFemjBD4yz18rP1stF5GEFiieJrIlAKnF+X5
Wes0GEujvoJh8cBnaTTdaf3radRII0HrB9c88HmhSlKIiMAhrt1hHdXK2Tze8JlMXFIKCSVve1HM
5hwTdBp3Bonh1ISrkGEv/Hz6JcV8AULQGGmnhpt41FCXkH9caDJgyVntjrhXPQ5Jwr/JOnJmnycy
RaIePR5goRB6iTDcJ6C7wq1/1CzmcknEgYX1dV6me7kiKye4ohbNjiUWD8uW8i1v6Q98tCaDLCDL
wWCdmhthHPpv2tRfedYKwyWBQ0DV4IoFt3gJXQsHAwkLwlCVjxoYQL4+QIaN/pkyKSzf7TEnMmUK
23nqp6L25dPWtCIU7wBfqFuLniB6xdMKnyKdVaMlTk1NgzpdMT7ucZ8K24xO4A5FcBNadXxkbEHR
BmUlr0nMOM8cF+n2ZiwIYsIxGGcJHmrri9VA352S+/EkFlyZ/wowWFw+ccJ04xhndcgBAtyf+CbD
kaHe0FyIdSCxmkHiAc2HErDsrr9rLD7skh5xQr7NuD6K6Ghb4f0gRxm1MAWlragAAXsnO0YYc9vp
xUgc4N7q7IH80i+WJExq4UrSfANOP5mhVrxKG3I+Z0kp37c0/dFmMc3eoY31E0Hd38UtCMXxVi3V
j8a95bI8r+nuhFN/d5ik/ftvxXt7MXlGvV480FJtiQC2M96lt68HER7z0AL5u8fd4+0CczwYWzzJ
CU01bN9gH2UWjRe8/QGCNxb41JZLLySNZ/HRPJfqlmvQehGgCexkSO0/doxYQ5gpSmXM2uowynxg
+PvJFH0B/BOl8TzhTXa/eV+sIjo1rBEGf6pewJoBOTNjMjlZx6vQHllUvCD5lJOzlCc8TFPysnQy
3QHA5AVMODXLO13hFeEeFc4iSO7m31pB8iyIe+/WwysfI5b1xCJtZQIf6FApCZaooP8UsZabfVgy
TTNB4i0JjoyGK1p5UogiQOnNsCBjomFkPb6ZWctZ1TUPh61kFK1AqngvTHOxluKui6vnkedfSgh8
2NL9dhegDEXkpwKNJgrj0ccMq/H4UofwMkUg+lOC6GugvUAE6nl+XfXj0xxumgFsmWdenNocF2O1
MZmNxOrifPSGNww8UUlJ5bC9qwudScdLqSSY7q7Di1oOsEhvkpmSXwfvCrU4c4DFnwIW1rH8VMvX
ZffxQW0C6fRTpdhvrUqlIh99YpfkSz7DNrroy5CX66BhVx1/kvgzZgUi+D4NijWW8tOP0BNJFefw
rK4385bFZITDSkI730vY5aLYTHFiB2TWr1V1viuPg6Z1YqGxVgCRfs9WK+08qapNeA9o+T6P0Poz
8i3dTKSkFgHoNLiIMJYNsUtSAU/zfJbxxMmDecYtxZ3xkciCAp5BD5QuA5BUgBJ7WnkFuR3sDQhb
QDR0ZPxFYiueMMDN36njWqGY3rj1kPxMsvAvfillXzccT4oAwu9qxqIxXC23v1Kzp54nAmVbfgYM
4BAYkm3SrfznpCo+lK7cH0N8SNQOjexsK9YyTQmEZTU+vECObo/BX/414s3ebmu5NotF42Z2A6eO
7CNIZmceFEBmSwkj3svTJ43ItUyIx5BcmrFh2jdBC1Oah04q8wPVukW1wxDr5WM1RSnqJb7iwmXJ
8HEOuZ5cVFwYMFy2Cm6eyCDHGzOL35XffCJrEPIqYDBsJup0clmsq20KwcGVZ5mEcsCvbdwDHomz
BXbKhrDACYPhQUHizqiLsTzaBGVxjUs+94/4fPTYddPxBXnPHtvPGlnV2xnl24LJyln7N8DnS9d5
ruodzLz6ggteIOSYJOPEhvHkyDiS3KVQ8i5HK7ADcuZUmHCGhl/th80Z0HUmB5rY/2iTgNBrz4/Y
2k91raGGcZxh2+7MB7HNQNxA288fi2b+YT1hodaQI6oWWaCrXuNJ2dEqysUTlemXiwmvv1EECuyA
uksh8dIdSG7G4wpmEY/PSfKXiMLqkjUyLH74ZI/l3MG3j3Mnte3MU9dM98kPEgikyN+kkiNTBZIQ
NkdWPlzsiCCfgKb+42qO07snYgcIwV5285UunJCy+kvJ7/0Bo3jubM3bb9iDZhgyNHlcLBJFH2F6
AFyccPx/NvsfW2yi+IyeYCYRup71kPFXLeiE1Wv+qXp6z1ZIwUErg88P9c6s9DYd7hm3vy8X8FMl
51CPqZ2p2hHdeAGPDDoAG/+wGRu+9OCiwpN4Uubvprw5N1m0tox2/hq1xp/H0eOAsAkxgkr+KBLm
3FcjrawAhLwcsNsdItMqknpDcXyAiQ3pZdy+iP0POZj24Keqw9/DLdHptQP6fx0zy5I678/L0ALs
AcJ0wqlwOKw72UfC345ssS7LWzeSRok1RMHyJlnLBFZMCX2p4oUwWbn490z44OSH/abhnmP8Fa4d
0GyEcG2ar2fVbv52vytpO35+vgOMY4/LVO0iffFxQrJPDgZWWcTc5rhc19rv36gzNjSyaxkAuM6D
9SDmgnwaXnRWb8wvOCt5fGueEFXhJ1Tf04Z+jpco11AEYZxSg6Aqz63B35NtAML202oEGaGtV6/z
b2jEOvjj0VHu+245eI1R1equrlj5YwBE7yaTsTfUAFMI3YY2iDpC8Av+0rStBnNbFPyWPuYwhF8n
2HZwL6IpxdPmfsQGa0d8vjHx1t+m+LWDfSE772Edqq03y0ua30ARalNy6n0s9ZZw+Db5pRnrdRUL
OE+0RAs98d5bvQgnmjzGetFZdSgGPUpHtby6Ux88xxdT3uEXLqlvrw8+LL2KPnqew28qd+5VleSQ
/Ptts67BCSNclx7sr8fR5ZIvUfmlpLmHyO9aNzQ05a6D9m1zFCcXk51uNGTm5zrXeP+v2+7UyULK
Hoph2ChPK/Zhv/rbGcUK0ffV3iK53B6BkaIHKkNe8GX4ievRZgmtQX3/jP/d8GXq32r/uIBnOPhA
z35HTFanlroQXnLrZ68cKt3lKt0/lNHnNkEsfLIldsCvs3Thrc4cufuvRv4+w+h0kc5PPPmKK/za
cjEwVMLnuDJpykh3r6nr41VztJgeY85sfz68hP6+RUvpDWJbLTGFlEJF4V9QCFFCpZfECDTOOSoq
TDaHt1vTuVOEVYnGl8p8SL/7gWhtIoECT7rdSZ4Q5iaBT+1j/uqFzTyWF/kA/SqsIibfXMgrqqKg
wo33RHtdPuM+IilPR1QVdeMemob1hy5zf7WVKNZ6Kfb0gJcXVRj81IvC8OB+LQ6RqHmNWSFvVkvC
4vepUTIZvKM2mgLuzLbHNgq/jMzPGkqjrZe8vzPS5y0Q4BRvzyC+hmkqq2t3+1sfCv/qBiX9rQy6
iQ0zoctphuaBv7ArQuPjN0pKBflBJVx3hpAeNq+Slx9Ltjib1O5YJKNS0F3yxUp66tWzxoV01Fle
BK6NQ4PiP8qlAJqjNeDiCnsVD3icytr+8MCjb+I+ujoE3wzuNRH7z6JLKqRPZ1vDp2bRBLzOSnlX
OAlSe6i5TuPTzG1O0w9hVYkl+f6OS8RbujZoWKAHg/8JvRygVNVzi1+E+2bzBKdlDH5HVxFHWcxt
B0dAjNA8X4XKJu3C1SFtcKpF9Vx65ULDUxBrAdZdWeKIw6CjovaenXZOUCpMlTaApartFos+IPC0
N+dvhTkNeUkeBnFImQE7Wtp4UI6Vg0/DRX5nNzROfPTNmZSfva7GXu4EuArg/8ksv7ETyLVPTtpH
RFFMd5EYzib+auqjRsztm8BuMph3WYNJAQZoAQ/48nFRvrRW4Ag2H5M2vq8K4sLK4jJMZyNAJV7u
zyuJ/lMRV8ekL0q4xmC4gN05f/A3Gcd4mbtXwo9HOKeco/4QusdbeZPB6bhVmhg8Q5Jxic0WHRwr
B7WVq8TgHZ8Hr0SzMvLmYF+fvxuTDE4NHmV+lyKijW/cQIYr1Qr4E/0UbGJ4D1WEBZWOq/cpQEKx
YjZov4bHuqSZIYHUw0aS+qPB43sFRHq0kygjgIxwbKgtRrFxo/I+uOv8vbVgRZY7lRCBHWpEkyvU
Q645fz0/fN0TWL580Pr4fCTYCfIb45aeHUhoUK+P3uX9Pl0aG0YyJuyp0sKRF7CrALqr0y4kVEhL
ltWuz57K4jhE71N5+Mft9ZB3fn0xs43aSEmdx4a7KyaCT+oaawuNfCwvwf250HiJfH9XR6wVSD/p
EAKvAqOKC9Q4BjNjNyahJG+JWCX/xgtr7xSHjKSTTWq/nniYZackONlGEX/aOCYYbaLhz1PNiPZo
xK5h6WuQArFpDBInRn+NPVmfdmKKV0Htuc0cv4V+VBQLdXa76hVFP7DOtYqCob0W/G7FX+UvOV9q
/9mkr67CFYday7BX2bxtxt1vXeRFQIHETOjba+aQuPZ4owPCDDks8U6twdz64bf+T2PG5LceaAQC
MFTf+mY9EWEcShc3hUjlAr4euuVUpnoF55yz2ikNUPcWLTdXWV8BR84HKluOy6k2+PIiSubjxYeB
Lx/eG8xaB8SLNFaJ6w/DKKUUlehF18B4FqAPMbIcosZZfDGWtpC3lhB567f8RtUWjPfCICPqgpK7
P3q8YAWofafFmx7UlyAiXu9qzwCA0qOPsQqLY4k2VvuLGcf71q7RaafbhzItulArqbWEuHr/LXpR
bEWeaIljnVD45oLrVCSJn7quYYsFQmIDeQtezDRGWirp+nglewgs/XCM/z6QtIV41XoRVrcDxTnX
eqSi3gPmZUAhpCV+G5VrzezdLT2zEmNjVscUToYkMYlGKcu/oD4ivJXNct5PVlhi6RDXl2qyeYyq
3EjKoJs9l8U5kRl9T73jT4oxBUnPh4fQLLra6xGkd6w86uIqRlzt0bxU41Gwp4jVXy5Fz8ojXuXU
N6UHN3Jtvzb1Cb3s4tVADQ+7WIXsflB2KFsZnNGnNyW3n0pP9iEdvdPL5ZrtNeMqCPvGyvuY3Z3N
pRPD8TI+pv6QIJurF8XUKO3CEv+mwZBN0uiXDCpvWZyCF81O6Vy7IQoJJvepAqyrw+n/o0ogLmjT
4K5VxOo/rg4qa4OJ6e2SX8clx4RD1mJ5iu5fn22RwL1AITQaCZxtfmjhhjCk/RIOMqtULYyRXXYd
T9jlyfSbZBuKyXc024/66HwdNOjv9OAiJ8+4gY9V6kO6veC/74JNkBMQNGdHVZoVEEeInimdIRcc
HdZJGDt8ZRHA/DFoclisOHtCL0elIEj75QJRTX5fyiocK0X8OFimoPvkOv58uBQVDep+YBjJYvq0
d6X+PvSJai5G5wDNZ/QUjTLtEv55irGzfDlXI64DvwntZkc6njm3NxCUIONVfk11AC3dg/ywDC67
aPLdNf6DRf1Nk6fJk6ZMliY9KD0E1u8lQ42paIh2BVLMcaEnEpy1GxqIgx6KtOgj2LWFBISS1kT/
5AAjwFv4N8i1FHfXMjOYEC2Rb9JwnSyPeZkQ37Xg7hiLWC7FRwy19RZvs1bekcDKZjGt9qW472cX
+m0LHZ5unZ0Lm2Sqcz0mKQ54HxsoYCfuUxuuJ2jnHP2rC5wxAFIzS2k33rB5yNx+0LalC8KW4oK8
BqD3UIIvCbIYdTuM7pX5gjIQ6vBZgmXlLsDRA5/G/IDCbUjnWD4ipSg4s3P++Rc4iJ72BiKve2t2
/WwIER0uBRSD0cTGcV+pgpYIcw3Mym1i8gjCgNU/dhkx61cqeye6tl2VZJhNFiaL9RjgXQr+ypAx
Jj6KVcCVfYncwoC7KGtRcbgT9EGTGm3BHkG4b1+al7prjYor4of2tUoOlEa79lQhWdmXFtMqIWEX
4zuoABPfiXyF5jxLBAJNHbAmF+v/Y4C7Qkvyoszm0DXZYJo6cegLv4gnq7uS5l+liQSZPUpGT0jq
gPihxOqC5TOoAE6Y7fD+uZLYU8AQ08eB5UCQWreFTcLGqyvlmAk+rA+QiHh15Qf//8X3hGSQR+e8
zWLDYV6MOMyMbigzujpc/X0SWRZux11IS8BJAx26YAna4Rgx0wZP5S8FNKnOsdNJnsPe1mIZfY9s
/Kvw7zRJyGIN7/8elvNuknFf8BymDvpC9VJJ3eFzcMR9CYSRR3mRjc/VNCmjFlN5kAEl6/e0ra1l
gjlaGY4ed1I+mG9nejlsKfnDksBK5/mI7Z8+m4nQ118MoTKsbhnriiciNiqeQeY1bYJq90eLBnuh
gk8saTNfiKi0d0sGEIWSszatSQyMvOH3Mmtify6vtQJP7A7pGCeDUYm4RMthxVjAxvu30a06jks7
fgH5tUGFWfs8PCOj3aWcGSp5Y6NaJtyWzuJ5YjSqkaxWUG9t/g/++UCQiqEoEj7f0+iD8+4WfVIx
9aAB6GvNIYwXyi938u0SQzfi0INEAOMeYjnnVykY8qNn0D6fPAL/LojHYkzDxn7zDBl890ufbUoh
Fe1IEJTGNWG9S5oNkemcgjl1PIqxLN02yXc7yJpeQnrIl5GaTb9IknzXBaFKsKpb9RsmML17dwIc
TTMs4KX3uDG4kb4pZ3x1JXmzJH4mSlApdn6wMD9XFCfBLVb/NkO1B/526mPeWhke4H1pe2LxkEfF
yqL0qrCkfgeZ43/HT5XeUcRjfdW15b3z1EqEYCW/29md4r/yHIlzRevgS4Ps77K47lebfhtZE+zE
IXnILxcyjv/oD6PMBX7MtTghMDr8eUqqNuj29LVf2UZPKzUcejhGHesSvHe/bgk6o6fzkBASkeWr
cBgN/f8hMTIUKemjv7RjVIT29oLTMKMP1y+DraihnTT8Gxa7gFDH6bFZf29+KK3D5v4iSyEoPz2b
rjBhA8C7pow/cfvSSMCOX2fmGf7h8ArxWO7a8rRs76rufXn8x+Ec9gqCLyVjSYGDl6jsyujXvu3L
c02JjOTIHVIjF+l3ckJPzCByLb84ct9wJdfKkk3GV3O9TAeoTTG3x/Iea3BHCJASlmFf+Oy823js
CQ7Mu/gXPktC/lUgT3/P9L7ihV844Rx2AMQhf446CnnDLByKnAb9A/xO8Yhangw9NAdTmK9tI9wF
gHWFTBamFPSXaPrpvh1B73kdpLmoXkTvLk1ac2b+LcUpVXUx/YSc2ghe8PcV/RPPAyR0CvkQHiAy
gmah86WiOuqhEc+n087kNAMJFzZ0i37ypobIlZQXctPnPu9i/HKbkdUkShnihP2p1kN7lyyBGSxQ
xkHloSwgK7h6LbC43bv5nn2FbKGySxhMLE1hElTuTrK+2gKbGk4URB9vvIq1UiXN7BIAxdxnwSIy
nlp14qLTKAG911cPo1oK3slfMXiiQgMjiK2rYwvUvVzME5E3d5YvWYDefdIgQ2/LFFEIAtTnIDfh
BkmBwCQCWnDehHjnb3C13Bw2qC8Obnh0NBXs7H4S5XuDiCK8z86usxAIOSMgAsSBjiX3QD4qut3t
eedTHbE42Ru5Vp7z+P/Du83qwiWj0ed8ZWb21GTuxHJ1QCEnDDLDjGJx6dOXYApzee2nMvZGPHIA
8MGeWZLTl68ox2MZjdwrVFO3NjK27ALaWVfxYN4KO1OrcWrkQodehBqcSf5rxhUgDG+odXf2yIe+
C+SwB5MQEgofBZE0FUiyGCMA7SZ11qR9hvn88Wj4NsHEqqa99voKTWygyrERZUQuEqTG431c7G2n
FYdzO94CidsM/VzkiAgyPOqJf8yCeTJZQbjonOE3knYePRl2qI1MXf8hBQkYSsNiQfwTwGJCeJJy
zw3ZlYLX17tHDWAdCVj1i9BirPae/U012TxvwyZKDmxWJ+XQ1eu7PNB/ciyOmBRbGtUbWLHbmver
bP+T+bHxTeYfmxiTujNo6rM/iEEFDwg53PDFwAVco3Loc5GmqTrO7RfGPPQMKzxgenzWYQXjN4GW
D9Sr8bCiTHGWbHeHaVHnBcGh/3mYr/R3FZZOOwck6YoEfZ7wG53mtDeNFhrASR/lqtAKVxSmbCGY
TXvuiVhqbXjMopKgCpZpoBMXUM5vcfJIt/2OijCPopzsYmOZ8w2G9KkN2ZzbuhqtipHsZBapqoVH
ujzLtzIb3WNBR8asWWFhfrgOSYcOXK4bO3CKxAigalF9gArx5I3pmUoGLC2dRcioyZZhWdlbe5+D
D3Md5t4iB8Ntkg5JdHpWhEiH9Z7imKBv7p82m8usByCk9n+lGPFHys0QFGDIIgdPFzh230+DYS1H
GNCibJDSOZCO+UooPKznAjme9ie6mncxcIbI6X1nyq2cvCY1Kz/8SEu6Huvydp6nOgJzyny2uDfk
UL5ktSTS2AGi5WbwLEr/k+iakKtDdaLSNNFFN6qfy+zzyktSbd1WB1MDbsEUFsIG1dugZysd4y7M
ckB+l/cTOG1mZzkhDgJ5BWdLVdMJ8nY54oRtQEMHoVnxlHsIXNtD6uthrvVGrMR2Un9IMWwq3vMT
NK1owy/ruNLJs8rBMOCOzeSsHR8QHp4TDVMnU53mPD8x8MMDt2f3JBwxVexTDToBRnT62PQGB+MC
WYE8IDcpCcnzf9/qsZQ8qNMi1HO448dXEpCKqInqGFff2Eam8wiNREj5YmFgNms0Dukr2ztCgiye
KwrBBw8amDfbWRd/mPzOi6sBtauo9HQq+9e7M5wuKs30ISQ5GvwBBuEf0V05de0ct4vgPHeMjGdl
9jtYHVJHgrbc4NFCWC4QCLgqseQRDITv8ZKCRF/i0P+OzZtsiMt661RAJHy01z8rj9Hk5OPxXMHx
3hIai2E1szcxT6eViR5wJ3QAaB7NauY9LxOLBeqDaCTzy3nTIo4O0KDYflZudipt67enz9t3UWZK
o1TFqBpbBcekTMnDZ7u0+YCWbxPyr+SKI+PZWPB2UWVEgi2fMMsX2dK6s8BygdKhPpBJhYL2csBJ
A+TpQUxwNUQRRm2BgoRnHz1Dxh4zhU7Nl8c+J1rfp2wYiEhxxYFiesTN/AzqDubnpNJMReauPNzM
N0Wx1YSQj8bI0SROLQMjqX+9lbSewbEOzgaIDyJhEHoGUskk78my/7dzZotiVjW/ZoFxAMwGc7GY
Q3iP41zp1TCoGQga3nH8rt2BWGuhNvMFy+DyHkwlstmG3rbQ1KaLjekNFl/bSX+0UhpUXvyF+5Dd
Hg4hpXH7LAW/2mY+EMw36ZNM8JLX29yOwXVkbmqlyw43lvVK4Ey8gqfGFv3+S1NWam23Uanjo69Q
ChWyU/FeDpP17FCbwbmg5CYGf5YoPRx8TEjzrSwWpShfHOPZkrihx1z86Ypuepg1ZrGser+Yh89o
urv/6mFL03Each/RLp2rJ6PAuIlEl+qsG3qsLL/8lZT1LEjBPHNTP9yx22RaWuB5Gcq2+PDBKVhH
6OP610CmedSIOQd9x45vXdN/WMOq8dpYNvqXXXosJuZAG1yhqCj3zsAAhmbE1kA5Spzbk5w36MYy
K0lhHxRfVECuEpeOtuCZwMFOJIJTi2YW9qQ/NX9N8CluLQW/duUWl+FYRBNhvsh3kZCFvKKuUdyG
mRglR2eJYYnDn3qcloHgO+L3G2B1OuH9l0cRuaop6bDoW4M4iHaJoJIPxMYSY4fACf4mcE69hoZ0
G5QrcW6QX01MIsM3/A3753jiaJc4XmsPxK+3Me9NFi7pMIVzExfv/ykFSOhgsC8S+OGXu1J83KZd
vx9h5C0iayMbZvDjDDU0z8ts1skYh1E9knF9S2nHEDY7ehXAjHvVrqZsHv628Zb1GlXhUseKKfHf
LR3K7Lthn78f5rWf9OTj3xkNru6xN5xxYhrFoRTriwLQ6Jv4XsvPKW5asMCQ5d8qKm0iwJA7J6H6
LaU1aEdAvSgbsd3eQck1hDQ//vntKJx2XtfpEXBBJu+bVEj+pCbTEt3V2Olgeaft+tLPWv6mka+M
W+lSYBqkB0jggoUx5gaoUK7v8PIXceIqAfGK8mdjo6nBOnHDlYRwaxs/hpbzZf1UpM/nHRZOBoxE
6Ks8fwfPCK+uYJ1OeAJJxIU5tYhxzUdbMtgacbrayqtGWsKLdmVnJBdQi0Q7ktju3+Ynleo5ezG2
Eb7y/kaC8UYnfMCdXHwA2HRpixt4RMfgL+iLyTDJ/Ss5+tbejxubBDm+P4oXyPfZcSwct05sz3IX
I8nd/URSC4A5U+wwaWh1MyV00T70gDjUBvPugTXZNYIMZzDsaXZ5+IvVVgXjns/z4rjXd2bmK/vc
iCePO068mqzR5llwbMVlbSTwiqDBgJmn4QRmkYKG9j13v8DVYz382aeLgUIWGheqUWp/kAx0p/u6
PIQNHBUddOzdxW3TvYTIVn1OcMkg+BkXkyD8ura5I4Pi6bYS2Krqrq192xdClLhsk7LLPzIh+neI
W/o2SiFznmrg3lvEUs/531RE6PpXkdCWEI9OO+vdwc/0lkCib+DHh0awtP3I0kfa8rYkqz0HWNhF
IHGhRK1V25j+u2paPlfixNAbjO49RmA9VJSwi0C5YfdfQUX0gJYF51PbRyc6eu+DW/xOcfmBmFtp
GBwG/UJgndJ+Cqa3eFx3Fu0EWZvDxKDgxZcgKJtnNc8M/M8SvgPahfxrXg4yd+4vfYXqoeC+ydYg
WbetgKNsEz512H00GjB9ytF5jJSbjCfv2vmyCtpw07UXVwFiPeFy3f4s7E8CyW61QKgyNgMNHy3O
X+NkCPa9HYyyGxJzA+CKZ2Um+txR0mpOSgMhtSKekZH6VTIWblWm5zk4SNH49GwaqNQBwXC/YIYO
awSSkXOr8S+mjir3mr7gO9FhX4IAA10dhULVdbXEJFFA+R+0m3RJeO2PKrfPPoz1GzTROTZFbewH
h+ArHnJlY7n7Dzs1gNVqZPRScVFGfuJ57aYUF2cAq5FOdvwwU49NBf8jUKVjfva9Uq7ryGF71Nel
M97hIjs7/TIcv+YFpfYJK4XfpVXD4mfciMgJunsKW1VwIJKB83kfLwTyCltr2iUfVXOHrywFCCvw
Sr0+42ILP7/ngFiB6C3s35g2vZLNDCX4rLob+1aUJ1eCyhj4VC9pxXjo3jWIJvK9zv5CnarNzEl7
IWQm8JAiG7TNz20hxdppXcJjXCixtEg3VD71ZmzluVc/9eLQHVVgfSv5P6QyuwdlmBoOAjRf1cOM
094QKyAc4p5pePvJgFpJbq+7a/ttaodYff3sRKzMIPk32GW405sDfs0/Dba5/uPl4CX/4oeEtkK2
h7gfFnR/W5l+qb790+54MMbvYRpGroa8Eq4DKyMJEHtmSDcGijWxOcnje6YuXeQS3Jl2eHJmzi0x
3Y42griOSLWp3ZVfb1o4OhLff0R6isCavDu9WsOUNrwrm7jkMs7vScdEPz/+2RO5FcFSe9LxSQHB
ld/ZT03Q5PoC7TpQAo8pRQ0eCGrAmzZVlmYAh2Ea3va8s1n1VIj/5153IhOtv7ZRZPYeZ4DiV/jN
vg35aQ/2FQrmqsQDXliSRVyzjs2gKctjHqGOTgok9wfNRCPmiqrJufVBFp1WFUrCrGpS3N3b5wSZ
n1WfkX/fg9MOrLLmpHsYBAdARaOLVYNl1aXAgL5D6QnlpPfVuYrjsPIjhS/OPL8/QvIicBhx/1da
X3n0iFKthqQEpKgv5g2TkGPjDH53gQSCjYlvWzsUgnejFxvgVTKNLj0ASQkc3bGBc60taCh3Yua8
lOqaijKYW9HwUl3znlpkpIiVqidbrOJY0/yQrSz+04BOqGMttiFIqCh7cicF3G4wjcPM6ftyRucb
jfw8dzNKWQru8/eRTwT6JceJjlvif0XTnT1359gRhiLJHMNK38mv0xg9Rc72TlopY0o/Bgng+AVN
P19U9MtBtqKRGhbXMlhhJJ660+d6poBPr8NwVUmjm2+AK13/3rICG6n+DG0QFf91gC3qzXoJpu0x
B8q6LIzF26Smq30AL48pY0pYq7io9xaYJeH9GQ37y2tIz0QEgTB6sm4k/A/Wd/hb/5BHMBWJQot8
2wFOzDRgZfXORBRU9tdPVkP7oFyU5Cg3RHQv+gVI0ckFjzD4/KjdmgFxL/vmeKWsnUZyhIjZOq6t
TnWKPXXkrIxRaq+zkB05+ezRvoF+DbQIgB6i8sjo8L8Aaqcp10pUdFcCsEbAmn932ASYEAND2ZBV
Clcc3v326lpjp0RIWOqfQNqp4UcYi20YTZFlrubEvCsWkikZ2Q2tN9BAsNBNB9TDRJgCNHetE/Nu
iOOCUqUfGBvqsL2qPKbewrJeD3VvZpjL4fkn5VKb7gFtAqKNDOUAC1wcNDIW4Vx7VAWnMQVPLOBJ
RzS59nna22gFL1zNZ10cswefd5eKfybyym7mM9RD2MsNxzGwZ4ZEDFKkPPCYQXTVjJfzMFJCEJGQ
3vLigWDL/x/ygD5LvqsPIGDeodZuEGb5Fw+MK0s0baqa8BQJpQt1L77IjfvSvNeM49McB6hlKON9
MEN0UeLrUHaPUlQWFICN3Sp/4rmRPMl2wZocXxGMqFIth3EjoC13vn62HzeuHcq5FTw+IkEYlVzd
oYQSo6O0QuTQxEWNkETcMAHjkIIfgt1O+ElQhqI+MkqOgfbrLpcuIaBN8kPSyxBO8ARcB8cp6XB1
WJQvd0hBCW5ZJF1ECwpvbctmsBbFJpFvD7AquIWdk6v7OWiafAQVUbyhVprgq0L7mP+r96ewX4cz
lbsQepyuHyMoZxQX3G18cuT86sxQkdPG2UfhHlEfJbZi3I/0Rr2ngSYgPCuM+R9sEkjf9gcjb3Bw
6SiKrRrkgr8cdGrN50svTgYfkZUk8Fu03SgR00xctSsohvaTGXnFtTm/IYLY8QeF4PJObcHh7zOx
KrymlnbCsduD+kFYlg0xFl7dnWGfe/nTgakqcd9bhKhGzf8e4LIZMvzoJcdy0a6/MJGeLPsJZuCM
HTqWnGsmVJMkHNsLfLMmZN6Hm+RPTMuzGYR8+VgPNnHO3qO6aizNMUf80OFjiDDePHFBtOlU8+BD
yPaE0wyaY+wZY7q88oOhGEoBiNSR7VNLt4d0ix+1hJ02h4eTUeF0JUr05yYVj8SZm0WWO3bemcMW
YBnWgXP4xJbItsXt+UJb/uJmNFVJ462gpXja2FotGx8DvheAn242FQPFfVepQF8wqEXoMAGRn2Vw
Z8Rz8nHhp2PNgtKkfljB2j5NU8IeAp1COOLXA+rAppBbMnjgq1anFDjfv18P4KGN/yumOA7wheQs
99MX67rDKZER6tMBowaDSm7T7/71W393pPDDVjw+fDR3UDiVnQMDjGCfIAYdOvVdB7/gBMDd1USl
JC03Ccj6EnQvtnInvfdRV4cXGBUro2Vefio1y8cZgJZ0CfN+HLB0aRe9VNNbqTzq+DQDuLKBs3Im
yEEwWUlSIzOwxXRtMPqphEvN5vTzvVelHHZFhrxf/TebhoWK/ZWs504lsc1tTscVohL1/zuBCHgZ
0MBvP0R3bVJTqjvMjjEC8ZmA1xuDTtbMphBMibOiCNz0in5cycxoaMBli4N+TpG8x8NX/F0XRBTT
vzF72fMUGf9PXJhOnS9xnsg7tU8sRT+ME0wcgrttW7JEmybP6d5+vkoo79rMFLwafcVnibVFBh4D
pBnwFyN+4RV8lsiF490a2xayx/ob44Y8L8Gad8MoOxL6pRsMhp52QUO/4GojQHc0tGssHXWvCHsy
C9TvIHXCIy7fQWrFTslXfUsSt6gGioV5qO/n4099cMYn/BGndT14VcragRE+RKs9yrCyJauWQLcm
RtddDYAmRJ1o8mlGHuheXHYtuang+Z0baZxvpg31b1TlPbnXJPyfkrxapTNl7dpodsnjRDWWS9Z5
16crY7G++b8JnIBe6Hd10A3JT4R8vW8kvVWwVauDf4CaEs4PhVjzS5IvHVSvmvvJ7nXNhxAj9eSo
N1opjf3JYt0+tFkEALno95gHr08e0rMzini7BfnTv0KjYwLROqV92B9gmSMqu7SSmu+KFxnNjq9D
mc8pxFn4QIAJGSjJEHKUxkdQSUY6Zeb6rRv1aIFOB5nqaSbSkxjPdnxsb22teMmSWbqDVWR6/z3k
VbsR/U7szTd0ICgA29ZPkq4mxCzrF4rhOWobPl5Oi766CwRlnqrF8MguiecWLAcMhPObcfYEX5CP
0KjMh+jlEA90EUZsC82OeECzfrhk7RQyVy/k14L1fawtEX/dxovIPTEDj73w0/Y35j8OA4f+dC/x
ugMyXHWEqhx4AOrXwIKS0sstusck5/U7Q2ooEMBzERRiLYB5LYXVPeCeK1oTdbf2uYcojrCXQO7P
lCy885ZQ9SqfQpNkVWJg5uUJ26EaJDDt38Ie8TyTMc2Fjkw27JPrK1Q1tQyZzQqnn7JPRaTKPJCa
DqYl9ghHBqqe6XTTJE6jW4DjyZKVFuL8OxSvReUnsYbT30/6uabDSzY0AXcO56S3BFLRDjmqh2+1
hRyuna7ktf8Zh/SIEtm2Qpxfjy2uIK8/q1f8JIVg8+q6xd31GuHGCGKEpGHj59Qoppnv0gqBrpwV
B1f83VJjlPFSU53POPmdV1TqkIoFilL7TXovajsEysvNIXuml7w4nBxOme6qBGXVnwPFCI6GHqaY
BfzQgfPGaV+lEvSGg2kebdC7GggJ0/0MSlEKQu/uCM3RU0rtbwI0YRyTe0F+sWFZwBlur6sonx8C
pPJtsFwSujLKsU2d1NAIUOMMhdImHu9g62zFh8Ln46XGKPzF71LnpgB9rjlnEriH0YICSnvP4I9j
HYUU0Pwy/nD9k+asCmvLBvUdbw7sItU2m1zdpPVm2KP5jfaJuTapu7Nj4Dra4qF+2+jUFUW68g0K
QqBltwuAgDMWkDrpTUbSFX6FNY/aJJlOBEanhfhTBC+mhL+gm7fWszIFkFi8iBjVpQPeABYn1vnX
zsjXbM0Dz9Vcvd14ZhkpTY3v7K/yyMqMmzUfhFrVPZRcDnTZyOEHtMO0kT9V0uHQrJzKwIm12350
Vdi0qXSiNO5A7eBl7wswD7zfjzv0NSq2ISKUS8HRNbjrQwKtVAMLOOH1eOz4o6t6aC8Sg+TDZSwR
lffyDt8hoRI0QQp46lvd9n6vKWShKdId4h/LG3GqVBgxpcTKa5RuMefNYuNqPLBcrv24K69qZ71k
qb2js0/aX/xTrWaSQaV7QwZYSxFQi5tHcw/Y1iI6NONG0+Vroxggj/R4XeEkqZS5XQQlggxYq6r8
ztC0TcktwfquhE0sLFCIAOWQd5x3RypWZwGfVZ3ubECPkDe2sHUTfWR376NiMRDH9SH5eQ58S7+G
mO6N19iiOx2HlYzmCAXCTRY0chHkJyDANrbYVPOw6Q89fG/KpgCuZ/NyxcYaIPkrST864CCc47lo
BqAk+2c2lnswmDnwe+mNHrTkxhFUFBaxk/ffSpjENy+AgKpV/f3gvse/5vQ40Gtu6N7hUmg2RbOg
qUogPgBFg65lkfiZEcQ0XAsbfzW9iIIbeQEXWkD91mxUXiKi5ulzItgvKmQ64LzrQATdwWw5a6pl
Tps3UkjyoIeYke8lypzKHFxF1xSGz8uAH+WZM/xyg+z/xQJB6lFzZn+unxrDidxbCmCe1jJaTm1h
5eNJB0esc9VZsUd7C6dB7pT0w+f6Xskj9oTk6nkHmnDn2r9YgBo9vccasZgirzs2UNDsEnykxS3w
jTXQDA/zMSn70JW3eSvbJOcU1G/uBa+B+Us9kYiyY57DIZIXCbYUxgqeGm25EnOD7ewuTIULNLBp
TT/ql2dIiqnmw0rhJlxbsbDTCHJHbPfIj/WLYOf6dv/uZ2iZkcIJCKqRL6rGAPjWIJ1D1k4EjOqA
TN8DPuyoX0HexK3Gn8BIo4eKtG0U9OqJzM6e5or+ePMbPMKhfhbd9iRFSyhpwLFpEQRsop+GXSBm
NwgKgip5JaSGIjAL4ftOPzr89OgMzRxy3S+4BaqtNc+6k9Avk6tiKefG1tcg2k/nJxDaqSsRx++W
O1sXNzJrydskQdCSQVGro7xi+Cjzc1R61nwDFl/2NRttOxRynH8xjAkRQ1mqcKL1jxuItoiH80Nl
ivncr3jIB75mBrGg11An4ipuAbukFiED4eUgxHwhLlTMEHUBUgi90bQbdoPGcjf4Kx1cBxbU90aX
hVBhJ5llVe+pwkUGIV+Lzj1rl3Sl4IYr1vYLP3jhUWmD0KR62KYodZhUr9J5twXPfa87/oLqUM6P
ZVBk7CT0QIGBUCqUO3ivnTzQ3RNU1cNhK++/MFqGXFQ29PlpY0uhbcPRncx4pN/LvtCeIffowrev
1dfqkHYcMZSvjK1V4w8bePbbggBulLkD2u4qmaYNecVIc3T1h7GcB1RAJdgboWz8LXhJdN0V5fEL
xZX2k2nNHYb6WZCr92UxdMxvoyDSLMoXb37Txh0B7FWUypxluE4ocb6ilVv5Q4/ZHBxmOrtdoQrs
+BPH+JnHwYFnhTivCEMRo2mckY6rWK6a7+OHFch67IVl8acaGtr/nHplJ+hrYExYTCG+hC1u7yD/
2w6EDPDaKrCf6PRXoR3sAWcvOeKi5IVE9rT7cxamCIe7uC1HsMTvnbq9M8CSFaQG6OxgIqfvb/p4
zu3z/0973NqIurXKFU7v7KWuibtl10PqdiySL1qvNC4Ab+jRVjRZqg4ZBlq1Rcuhq6rd8PMuExB9
/uMym+aFJN0uitKfj6XsiArua0N7C03xPpTTfFdMaO2r0fw/RXmQebN4FiKCRPbADJWz1xrIs8wW
Bs2Z90mYp/jvRaA0EV1cPUTh+ztJp5zHtSpRJbUdK72kjRD7iOFQz1JSyB0PKTrsQSDaT8NPGZxX
XzeFdpRw2XktZUlp7gr30nfWZsvndi3HyM2eqD1BPhyWV07oTcigaZ8hwoywl2mYe3/K7NSBsP0E
rLxDYcH+1ixajLIjzniXhuy48DT1tiACNrZsJEOyFkWIVpbCI4COUhCARXeaq3GuHuYJEEtn5H+P
xp0WRRZucbvqyQFIOEjKGHQRgnqmDhP9SBTECwPgJX4rqLBB331sPZ0NNnVymqZ4c9pNEmYwRCej
2YFAGjQNf9ZvdyQ2xjdUCmwCWds44q9qIYVG+hbnh2YP8fOV+QCHKTjdFMVKFfLUltPw6n9ulRV6
LkrtVhRPNoU1cjp13n6mWM39Nw+ZhxbP0PCbHJhzYmcQufEHCUenZ3WkM/QJipPz/IzcNXXxGRtd
O1RCXJH+rqWjn8dOfBJXnq7Hu7y5xVfjHdntC0vNy04w+cP+YhG2oEFjGmDkLhBzkPgiX+i2+KCv
QGJLqxrzCfdGM19/HCex2bD0BxKnMj9O4Ke/VsOCxEX3xPVX4WBNa3UR94AgN1kJg4p88lzE6xbj
vpPX5m3WRpnGgOahra4TaQ2U4HM0NzFi9dgIr1+izvileDyaC3765tPe4ZWurCCeUeKXwAt88j3O
EHlEdpDSgWCz1Qine7QPNMRoEyfYMmYLkFZeTC2FhZ+o4MfheY4vRn6pSWPiWP0JCwJoiucrenA1
cYDlDTi4s5ejOmL6iXeJN7162f3w6t8i4I2KRCi74GKm1/uHYo4Kazij87o9/q3+GuJK+BWnU5/2
e7ypAhJze/GtYypwC2eXqt0LoFcaLqt+zZpHCYF9elBuipnx9D+y+fEHpduwyFYTP61dcFFvpe6a
ikHSP2ixG+xYNMoeCsCSVHC0ulCHINJ+vj2hvbzzhe0h0x694+qOLKa4erCvxtELOlsXhwj+y7pK
qZ4OteYIYV+oFoJp8+u+7nJJPWezTVD8iQjFG8wFrfqGo88KjkDjdzYIr0CDUKgVrbZSsTOSvwxW
JGkCe+iiIDjKg27QGNi7OvxNrAo6CLWJuWgqeKqnUT3Ch8KutdxHHAjHxiTUneKre8OS97+6xor/
8ryjupxlPmNTMhxKvfnerBOr3z8u9WXSQ2d+B+a4kJrnY1K66bKLDK1Yt4276ieJIc34/jx8s9mh
RAeodwUVvJUPGW+TiJ4UbZhK6E/S8PuUnk2hf7rJcBAjD4uVtykH/UoLYHAWlBaZrXzo3c8UEzrh
AOZPzVo9rC/z3bWdWkR1uYdA/j4Q9dLEyNMKI3b6mMuQnVUVBBG2rz95CnDpaiLFw8ql+RS0haVj
cY5F6M/FqHVAKizC184zCaStXPpNYSHBy8pDX4dcJOXvkgfGak6W+jgIkVhoCJ5tWhIF1gRl1esC
NHLiNXMRyrx3PZ4R9ENM/EAEJ8fC2EBCpSp2jjni0yH3u1/PzDLO2oj1Fuh7pFlgtbZxGWFuG0fK
HTWW5tFZQ/KDsNLS28J6w3JS3p1c8XcGpf41pcwzPXLHPOFsuLHkosabGAPJ/S20DrAP0UzfkRkW
IT+R6Rh9AHXnyPpD3cmqwzQ4DuIcQnMiOYCkvr7WXjKfz1i4BRKdyFXZOO/PiKUbNpc3Nms86Vn4
ptSJdKYvSKQ29J4MntFGGl0JjfV4oUwyEHtlxpEfeliZkCJvDnEL1nTwDnM8yd6B+qnB0k7j3MTv
Phamr9UhgbMRLvkAV0yv7EsF9MSzkLIU6DkqaXFLeKVfArV9Eq6EFpyZE9X2zNfhHVSYzLMPj2+A
ex0ZNImEqUQMfO1mgEHQiuCriX3Dkbvj/Q3VmBrAy4+zJy+lmk5IIbJJKbKmmWBOd7LhZFPR6kWZ
ZHu0Z3uZpG7lxDXbVEcfSQnkkI/s3RhozAw0Fb70YVz85IRmdhpFOISZWigGyg+eFPj3a10cxUQk
c9REmPCUX1LSzfnkivvIkqpMR/ofiLy1Hoax/9vgZQrkSJ9tg1qv7ulpUOo5KzDhR1yEd5zANlb1
9c1KCqXIDXAjEIzdws5GSFytSxz0YrEEgQFtfk4u09SenD2RqM309hjkEfZfsCCh3uDVsyNrG+lQ
XvF+h5t8vt+NQmPnExFQ7PCvWRGyLOiQxZtjypWc7xKUGMf3ILFH9T9S3c4M3nFnHzOJAdZL9/Si
VJoj22PvRU9VhytThavMLFFSAGq5/6newsYr+F/7q9cw+NIoXOuyMjaNSXhpd9j0mEKQ5PsnA2K7
hqJh5Q3E4EAeInOO/866ysZtHS+LpLJRF7kphA2drIiZyifdtHo9isk5nIeZnJnucXvDQoUMUhbw
LwnKcPBq4Lkv6QZgGktGnh12nBA2yuN1QroHzNPjxGYY79nyzclBy0XX9o3qYFBdr3kzTjEXw8r6
HOtZd6lv0fhoNc39b6pP5wbnn0hMercgzeKskE1itfSi5/Qck1BntNAYKspKfS1XIfntPEHdRlFo
FviUb/TMIwaWlh+t0RGqc3NcId7yrb5Z63CPqPTGfNMkNT9qATi0YyB5D+uVuttijSRzGCCuFsbS
I1S49SBBV6YcyieGMLbWopooeMS9lmsozr/I6QiX/kmHxTp0UNj5Ayw/KIpsCzC3flXQA+XdUXMv
xj6TYmvLM6DZM2ZAbwPE3pD3rpL1CDJpzmKOfWvEiEDokl171fGxeUT5cGfPMna4ebN2hMX7HHMU
IuG201y0yfGhBWPXQq4w7oXBk35ROnlFvzSOOjZi5+2Bx83BuTRxUIYMPSMB0sq2azC6y8r1P7Hd
vfVMlpeilf0vA6cHLTN28aTnduRU/IzERFk3o/xoc7FLYkjyU1xfbfCzzgVUHV6s4POJCyqT/LX0
amBC+VhF3zcJQPPR/mtZR+P8N2iAn+k6pmOnP29SyN5VFQ0es1rF1RZud78FvqGafPxSWgeyhK2m
znl6FvHLLHtRloYtICq3Qko2zaS5TJt+aNMJvGA26f5WpwEgGB3Ms2dHtnULttDx9nYZU5WvyD+m
dx9EKObz6/8oNhPSgytA/lh87f4BBlLr9aoQBFeoqdfkiUxqa+J6hjV7wQqKllz0u8frPhMcJgQo
5RsdiCFn+gyLQMk9MAPjl+wQIit+LsCqJTJPjw1Y+iePPd7sIDjGTm8BiyyJ8Zafwi1rmSNBGYqE
syYqDpzwCwLf/6JzCEPpvzrgkI3i/yw+mlFcqV1cxAn37rQf7BdLml94Ad6RIGqYGgfpGOltTTzn
ZMXlK7YZNMwFCqi0z1n7emRxE78rHZ4SdWj4834GGYvKVNeBr8/12gnpng0ApUZYcro+BLPMFJU0
qnKh5B+LX5EswIJ4LToCHyAByVp2azTViTj/Zs7b1P9h/vadPwhCf9MLPIVgwNpwCF5PLWVVYzgn
GMSK9y/cKVNiJUz8VHdZBI5qH9wqDeGsbxGN6nEuHbxUrqvgiLkLv5Pikd+Eb2DFcmY7+kioNEwV
V48Rt5K0Rn/1PcVt7br45olCQ/JA/UpzY/xAOgMir41OUxs4hzcVSqQ9yLe2UFzvAAth+D5/EyQL
xwAM+x1PMI3Bs29aKaJImxGgfYmsgYMzM+Il8nwIR0oUjjItBSHXchjyeJ/rf1MzEhgTkizTDxSM
562LGfgbgcfl1T+loGpmk/FWitLSg287wUlXR8auDTwS29JmtXERTNtE8rvxBTXwcbnfvgWZjBZA
q2sfRtPGgu1DqVLHYQKNYJwdWi+5tSsE2tINKQ4eeVrGwsWiVgAMrH2By2QTNPj5B3R/3mnqglhW
S4YoZhCdcWyYMxrTRAdHwJ631BplU9jwJgPwuPdeUzkQBWFs6dUXj0W3xtlZMJmtGl4ill5D0TX/
8BVt18rhj4heSleDAl89F8l5/d08y8nq6E/BTx06OdhDS7Szh6HX3qL1EvybzSi4oJKBSEWLA7zI
NfcbGM5DfUsIbDQvdalfntvgj4Sd1hy05q34vg8IH1nUfZ5wypUpss/rLqEZ/7phGuVaY+NcFbE3
3TsbUH+nSpgSKicBTTb9bcGEeP5+K5OMF79VzBXqlp6XlPKacyDQb0j6l5tObJ1GogdBt2yyE/Rl
h0EB3Ij/S320lmofGGKD6AfN/I8eEqBxgCC++ACxON0b7AdgC/HgA6wtj4UQDKNDnevc3zZN99J+
EkfO9SJsCG2i6FaWmHf4XYM4jkV3y8w9e7sMGxTFkDjIkybSJaAKtHQLqgScHokxybvIshuFfIrL
o9L/ofyzMYx/oO4Z4MiwVe4dkH5UuB9wCPnM5cYGNZx8cYBLMXKebFnLnAR6BuhEKefHY8neTdSB
2tJeoDnrSdbKftLiYY1T8TyWUH/XY6IA7PKkywt8+Krs8n4uty2rbo/FhUGrB/epKCvTvZY9orIc
Pw9rDHSFi0mYvo/Waz2MlOBYhMtkaix6eU8b0INmpZUpgBoL1hx6tVkVaDDPRMOG3wjin7gCKkVW
anN9GENhOnBTCIhB8iRA94cuEPaJBzHe9I3XaA57koXN1kNw6LC1AFXhp1wSjrKT3+uvJVj0SKhT
37Tcz+ac+GacBqJJqv/lEgxy7h0vDutdQ1kk9KmCcuVXcAGE9NzsgmutCz6MU7RITYp4ynZE38Rg
Mnd4F8E2eHPPrzbAgSe3GUNCv7Tm5lRPesbJdElAnW8aBQYV2Zt1ZCjsOX/BfbgXvRi8EC1320AD
b2A2D5llGZqy3Nq1tcQSLcJixkYpf2g3V90TsU7Sb14KT+I5Lvq4qgRYP8cqgHhJvjxJkuRgYUUF
f2aPcJ4uw3D0GHtY2/OZksGZ36QLZvDVi2ZQ8D5eX0K5DQ1GixGx/2m/QE2g2U3E/E0ZDsecO3Dr
2hlMIkWI+pRy90zluh0OpwIsYUUIDqvGFIwB+OQv0m3YRXMkxZW8M/gpN8BVZksDKTMe5HJy5uv5
kHKSHUhWCllcIhifvj5iuHwNmq9TMJjt+/aQwFIPR2NxsYFeQUjgManCtXngVmr08BDhhzKDYaSd
bmVaVJW2AbH0j4Lex1ZSD1UvNw3R3LttMBP57kW2GNeRQVhBnKH8tg32pIGwXI5wOUw8LbXYYi+j
hsZ0NKy3dto1ZgREyNxv6JoSsTDRa89mo4IxIu8kxnepyMvc9ppO1Yk5qf6FhEz5yHhO8ZFkMedZ
rJ0UGlVM0/L2Ah9HUrFpmmNlJ7ZVsOp2x4bpW8sxZmOY/Qoshrye3tubE5hCgTPEzG/G5Nox8rEQ
2/j95sc77iHAQSqIorv58j65JzdnpsNsuBdl2t5VcZwKmX48A2vJ6cUrL4zI+UKsjEISE4aGtacW
Il/CeLDurfLaifa3s3+7DqThk6xkuSDTi2cVt+UekIAmk1+sZy79YnffTyxlGcdH1z9TX9YwvW0z
PHTN8CdWY/E3haN6Q6GIp8QW4RPmTa7oXPbIAVPOmU69FMUqWpqTUYoQ86W814+nfgMGCjCCDP/1
QyB+zrvJ+7gYKlqaTyf+4n0FqUOYIZJWqM3fgpja7TL9OnTNUfIYp3Uxj2oa3QpMUYXWB6YYqDxD
dNpue7M+op+NpTOO1fYgXXiOdkiVuvnGHJHDPAdZDEmGb5pkcBNGZF1W43+BpB796bUGBtXmITrG
Ru3EoKWkTIfBDg/ev+/VlIKoAbGpTONDw2CZWaYIQTow0ddlIGrRDwzEfNkkrxUmvT2QED9ASqXt
hLTTUxoh5sHnIucigyQY4ebkWQvpd4fkIwBEu39yVdmQMDj5xEGI8xHOnDBiryJ0qBAPx3MHw9vg
NeFpo4693RSeoEfTcLxKyllRxZpxBNaijsxfRlSqOjEuS5+v3L1ThIU+Adc7q4d74Gyoa1kw9Hro
L5Y2HiEp0/X/fWN7yWA1m2iKU0XvrSpBzFIp0Mq7lPHWB1RJkNdJwJ+mvSaja1koFtyH424Q9Roj
sD78wPFmUbr17cZe4fiQJ1/7Ub1vdsvENBWkZUaaXFG+OsrfaYzlPNf2cH8G42jFUwmh9p7d1V8t
dFmsO0TOt9IzlcBBsr431EoSKQi9hQv8drZIaw3FaD+7THCdJK3Cew2AMin+WYijCVUVmEAPEhhz
8MmFKmmhWunUH43A2fRFfoA7TRRfT/iwKZsh8rxTRIHyq4uq+EzQXPkOY2s+C/OPg8dzO2eNOGHc
3JQcdt07vHkfMlApfwsvj76Fl4b/U4XL2CnZKNZpx6DQcykMOWEKNbNFYrFMFPBTr6t/VA1hamzf
5+tbJA0XL9+aBIiiIw299Ne4fkbSTfcheEqjcLbzBBUjHRKGHc8B3DFfrRUDfMhe6tG+cjg8624q
vnhr/uGkBbWkQUVBKleGNUlHTcs0VT/OOaGWD2VgGnt/GeB3AcG8dxug0Bzi1ei69x7xaLg5ULQl
a9LSE5+ZJuf7mSILx3UNwWj1jtk86Fvs7WlI8zChpvw1xBNqUbKQJK0NadMZWmkBHfGCX4IPb9Kr
UIyFGtsxDbuwunPwS81cpRPJNZPHYVH3fJWTv2gRf+Wq84Qb588ShhtlVSQarAS+Es0+qcsp4L12
v0r+OjDmkDdd/mEyfpI15HG5gyrW5OV8Et9VuZdLNbbz57aFUB4Z1Gi6vE6Ghkm38PKMLoCRAFg0
75eQgxbr5vwXNybIwCxyYqpH4owxEFybPqKd/u2SuN/phbfHLGaJOSFzuaadLNOQxRR2/9LDOc7m
wVxQfD+Sr6zHStQ1aHOfc28h+zOX3mS/nuA08rTQcBHS8Vs2EKcLq+I3Fb3ugU0KiA9TpJRfSBVy
xSl4Bomf/xX0Gvm3zBBkLQ8HzofYOgDq8Ysg6kQCvyuqCZH3Oc1mPpVF49dwYqyCyPwOsGyegNcE
gxsQfcl80spSLj9f+HFqUPxHL7jQcRtmU+iiOH6cyqtN84DLPuCfAtnoL1HaO8FUz1PpuBc7S9W1
SwgI7yPclysaGo89lyv1/auQTDkKI9v3xpu9WzjuWeapinrtd3hfpk1P9eV7mJswL72hYBKwIcb5
+dyfu84eRpPizdq/wkcmIhhLD1z3l8lzL7lexx9dB1RFkH/FQiMEJCQ7Ys3mcD/s4ONUJi2dlvq6
NgaaI87/fKmU88nK/LItSDvSu7wnDGGsP/7LZYYiMbbp4G2HAD8h5yOG1eEYg0aEwGL+YbCt6Z/z
pneIJkhoABJyVWdLw7iJbWmEUhISFUmyIn52muYcfan8McroJCaccPDz2ISHSoH9DTEpuz43mb3G
Rgywf2v3cWn9n7c5MZ5MGGdYfiQPrpvd0Jw944aBLOE2/qKq+0vVoSTubua6cy/NxxoErN0lap1E
W+crqnxNExqc1Ez/fk1yHgIHl6h2Tw8cbllF9s7IXi4NVcEA4uODG8/cr+tDdBBceHzayJsBSz/n
K2QuxDQrWABvhSh2eRTNzu8NOLSEs/eQFdMB22vS/mtMGZBUUXC4cBkJ2LRCTDAmBS6V7OzIdhS6
RmQWPt51JNJSk10M/39E0qjfp/SnKVVQqZ/fYHxSqrEWPV7cpRGNltj8ZHt+M4Hz4tbagQrh42Fz
KxN6a476N5208hOJE/2BSAvdaFpJDHQmBmkkT+StLvF4wcRT+U/m0COwE9VoarJYzgIF8vxQsvix
cLz1S8lNQKGRIIii3FCzvFoUblXjbc1+JGF/elb/FzxW3iDM4AeiBTIGmSlfAITxrtGDVmUlIXTk
jgUBEIvvhI0ehow6bjcVsphYz6M63n3nFbmvSm9ToxKqdMy669tKaWFpSeJ01+xMTFh61bTsLvXZ
efo6+Q2CbgYJ+SdtpNPxsAhW2MMTzG1AR2EjMDaiKqEdviBTKmxZDlXKjYTwUQg1BTSm7vIgHKm0
xBZhUyE5lbQ4s6ZCbPA3qrDJLurDwv2umYhe7nRbK2mteTxGLFrrQFbxPZHh4U/BEf1xn+BGhTLG
2/92N0pEEz/E1g5V7cnRTYgYZPId83CAC3M1aHXC5npQGRdVmcwXyewLcfvhYkiyOl3o1NQL7JjB
wKlHFSqI3cZRLDbTU+hQEaAhAfaq/GfRbM1c20sb/NDpZ/jJchqJpZQ3NFmc2a141bIAwFUgkyuA
PcQ6eVs+aXoyCZMvqSGJCsecT7bYILhkmCrcXGWSLDmfbPNRIAmlrGz3U2d46wqAlPENAaHWIVYo
Dw6XuuLMXYZ1yznAdvp03niS9bGh+UVfzAb7Aw2RcD/O6FaA3knTz+FYE+L+mU261dL998VjI99S
7pitefmY0r0TD7PYU82cIn1pP4z/PY+KCzqQ4zBRPbdlEqrzklmUcOi6NBJkCIlsJSmExGMsRLo6
xM0UXDTnWo3+8jCR3tP1l0LnDUgBNW/i9bdVvI9oPc6zi/1LdtfTcDMDnZsPNR8gyRBRvmB7Mt3K
OdN/FBxJRhEr58MhzA20vF0tyQkVw5PFJUqFc6K+enhqLAaxizglU3rBG/nhR2kS1m5vWeVo1hv1
NvNbn8eO8mvz9E6dVt2a+v/VJXANhbbYXAWcK9LJ3V9cee3hzkgqGaWXsQ6h/xBIL23pFMCmUU88
sWTLlq6Hwqdfj+2GXJ3E5qc8X5jMIITlg/tNicLJx9hulyRCBR6S6DdeuE+9Db09vguTwSWjbH3q
21fMjdurINmXNi/osmgaMpR6aFZ7wKg+ROgoj9oTpDsJ2qtR8sbeqjKSL/L4lI8oVKUYmWoJM/8R
Tta+SQfXwYq0wTk60X7rbbjbZCb5HTs4NsosmWUYe9yyp8W26QH1akdG6gszwvvUjKytaRc72G/7
3ntl5/cqhj5CyF9kAKcTtGihAgKf+hyxGeG+y1NaenRJgSyYphcRsijTj5hZPWsdCS+KR1zConW6
czyBvI5/wxDeHGGqg0JVTStLj32F3Ag146lUXXfzOywru4hYdfbpU7Tq49RB1vOth6VsArWEwqhG
SvpKt94wq2qPJUNYgQfn6WFJLA4gpz730ouONwyIrL0fj8kaVZoZ7S9/BylZCJLchtxvHJw13ael
O8dju2ne+Clh7s8qhEEGbQnmamAXP4+VpmoQ/GUt3eTSdVqRBvWh5GkQlbwbNmm7d9HF+OGCfrq6
K6Ca7XeV0+ASbCiM8UK6z6dQgLp4t9uPRnszgWgi6awTRhbatZ25J9otB1dFDMrgPOa0EV3oIMsb
GXGQkMSW73fvrvdOD7gRmUIvcQoPbPvq04gihE2vmzY99/jtVYSs975WOHP48e+1m82cTvb5yP6L
9I8An+Y3Ovk0dShStp5u59OMwDG90i1IjJ4dKVr2dH6pLaYglDa8G21m5E9Ubvc639RxJsNXOuHX
es4zEn5EIjM5ljzo5tQWJrzZ9m1CyMAr3jWV1VZjAOGoU89xPF3yd3JGzgLvu0W8yrQLjNTIwJYR
Vk1uGESkoEFR3tbxyyCt40K2/Vs1SabRwzOnpTp5ByTdx2vKRJtdveo9hLa+yh/DGdjOtKSZOIvR
IZW81tztNQtg/Afz1hIQLnuru+j3px5us75BU9adprIW/NV0rULDD0d/93J+IRkwk4Yfpmefi7RV
XLyvJ+E+w7sGwyPCy5fbiX85XDMxeXM3nshGeT8kp/2ul2ndmxoYuFeEwLZPmMSiGr5ZvdmESq1f
OP5BuQ+TKXhyBbTd4vVJJr2DoZAwQGbH1CCZzO9HHXB7gVu3Fx5YqXXD7YDNfTfrt3GkCURmIEb2
s5sJz1K/2gSEUIat9Q+0NvXBcqkdUY/jmg4PAAPUKso2E6gHrlguE8CrDCE9x760CMJensODq6zB
kyi8oazVAbjH1LAFp8idtAOYELspquiEFxd72OzhgfiGuy9NhzMVVI8/Ou2QjsO4+4WgYd29oXXl
hXFYcnzif6z5w7Q/IyIAlURYlatNkIi6ZuFPZvgF2KkWZ7lH8tg2KVto9o2BTDICkB7CH0JSiQI4
1xSKHvsW8WLv/GjzXOC27WKuNuxc8AyrHCYZDg65ntVEf2otqnx6o1ma8+Q/XA0k5tzNiKptrZT7
PHeeWrJ80ylnj2Y/d5V9t9JfBoPsTnxam/G6wCqOZ+Oa54RwkyAePNs3cw3wsi+iuRCjrA1CY3YI
ATM1/0NrnnmNcBUkJ9kEcOUsBfGFS/f+71ftZQAWJZ7DY9fodiOzxOmlM5Bnd+8oJvn8AgiZuSgz
zTkTYfyGhQbfUAHka0SCFVtuFMHrK4ZAz0ialNLnDlNS6dXV11Vkirsqd2+PIB+NZ0kwkiz4W5bu
yjRDpEvpR6Kip05BB20I4m8GRR7IttV32Uq9uRzlJVX+HcojhujOSPE3oF87P+uvD6KLo46FJf27
0GZjN4hMvjQss7y+Vv/SmF2v0GJlIocdrkPpT581MBxoSwWXrtxBiqqc2UzkjbTwdpa0QP47Yv6A
gN0BiXeyMZb5bx9QJvZgE/SXgFqR5RNHJSWcWtx+1PcwDS8SzkPijNv6GCV6HpnW9gQSuCLq8Z9y
F5HIAN0wS78Ap+ddvugqDPL+DeaP8HvphBcaxtJpOR5Mi6vqWKGjUY8wyP9iTghpKcqo7pPOLLxz
jnPdhBcGscUBqUSfTC5ERBXYpH2Vr17nWwXde3GQjiAMYRPJWJ++TEzoAUsMP+QSOcWJ6tyeGC2w
mUT/fQ6WQrFibSgiwkVKUs3yUrCkEkor4/cDiYuhbtFWKCxAa7etUlFO3Ty5IW8mJkhKwdSBVIII
wbx/oy0aqSKI/Ft9gr+pQIlEu21EQIfTSZ6fpoYCDW1NL4msnBc8abcyW69tx1+WA0hXUXO+r5Sq
2a7Sfjdotl95k0lMqHY2uDAXr6GBqTQRQi8TCcsomb8hKoQs08dlm8qxx5oLAqZdsplQr9a0OR2J
7bStjmxMu9cbKm45ipVN474IcZ+LPE6nmfXNrYt1kVSIM5P9ZIa6hbiHnFbg48hM/H6/tlJG6NRH
f0O7YVI3nz5S2zIUmUdHiUEit8AQMDvEkAXIL+DfMvEf8O8ZhhDFBXp3VNP6e9JTHFL1hL062vP0
+oqvpvSWySSACcCDX+ALQRROTMLKlTFQxhEeepLOq7Lg4Xb+KCd/UaM9bYTJ+cQgZAPLbedWbLez
5revIORX7Q2X0PQyCpRRuTz/wI/gA6QTIHxolnoVQk8WemaXEz2FfUoqhnCapaRo77LKIRww1HJ4
t9+k9G4Cyao26VRJF2jmYT0qHldl7jJOvbzeEJb9ETdR7WMTCzi0dqUmcUcSmLiJn2p49fERhHfq
ggJ6EMI4lShaloNf/neu9WlqdbHAZCd1AenbUUROivXzN/5eWvQp59bScWiN4Ao4mTKQMfqWJlvB
v89nnNt5G2kWSlg+JpDYmLAsTuJFJun0eqBG52Ia8TJtMCEHpqq53e54MkHdGvcJPdoOlhRVosU7
iI+oxxZw+/MwFGVb7R/c5lgaPyIIYovnn3SF1hhV9YKPJjEL5G6aLiimJBLE3p6+pAyGF2j6XJnY
I5RS0vbOEEzHpzM6Afjp8REQHRdhJiNW1IQOyo3miktLksqDMYVIfPeIu1Xcw06608ccj10LEvR0
f37la6MrH3jpAAAaOpZ5PNOt76eyLJLJ0BY8Q/BODW61OfP2cHB9sTZsCt5aEZeUl/6gnT+RleDW
waDKnhtrA0H8lMiRXbvWUamOzozla3f2/GqDFnkNMQ+RCEJcvE6gT3UgttwXDsO6WthTwIJHbkrx
adqpPtsVc6OQXNV7OfZGbA7iN7RVburicz98+FRw8euYbz329Y4GU11h+cSJ2XHtcib2EknYfuac
s+FFLDc4Sx+2Mde1ODFQT4EtxjuNaaMHSVR5vUk11mwrn12plVhA8M6UUk5H7sApy5g2masMtBLU
u3XBspVnz0f1XN/IczXo8TsgqqWKotGhClHbPOBamJbjB2aGDM7+ogNVTSFfmDz+QwmkrOYeuXs1
e+h4c9qbO02tjdgaqfuAsN7PhM2y3lak02REc49hxo8sy+8jvA2IGP9DB+3ybdbBhN2IlHGBqxN2
vodJYmSQC9eyJUfIc1WP0q7/8BkXpvY7c92XRzFTtXH6CBAQ2lAVIzirvYLJDkqjavwAPywk7ckB
rSZ35FtRz9+GNyux+Yxn0SolmSlzteFDxLCgQ+noNawqLibrJeAaT+oS8Z42FTm6UKO/g897Xi9S
H2urCV4LVjJY8GDqrq4ThPIkRujOe3D9iS9c/uvEHiGhO8T/Feq0RkusyuH1b54wZiw4N+HdW5B5
64u0QvxultPVLizD5geMwKc12SFVfR/Xma3W9CxDGLndnmEKWEzx0+/RNZiqJ45rn2KpnH3Oa8hh
SNQZ0G/1BbG0bU/v3CFLh73ELgnZGIMIQLAZBCDcGyxHtQjk38nHB1Htavx0Z0FbBMrKn5NjVlK8
7vHNhjSeo43PRvGBWeHJB0rNaa3uYHR/5+Rz22Hv78OfHRJ4qlT6whQyEeG5gvwNP2vnzsZYJ0IF
HEO4BPr1p7oJQCdPNJy6s7mXmzvkXYKGRVPjmnjkz9J9hHRVL5rxk3KrY834mnuI7WKgnVNuBHcX
UZd8XQ/f11U4H6z/b0+BE9mPcD4HYYvSKmwRmMbod5I5tJZi7Gv6mvMdyR3Wo9q6p8X42crozjnX
I+fhCmTKVUeB3MAENVZoUGePq3G4N0SzOTJ5Q2KC2BpGEVIWMNTqI5iNhPb62pVrhZ11xigZOvj7
1Hld8f7btVetGsQrtAAby1p6TC3ZYrYwKxOWTtEuRc70oX9c8bZfKdKLMxUnoeQPVdIGhhuSqF9v
kwpbvkMEkvi5sQhKkaS3gs+cPjCZx1JxLBFpWt4OMzLdirCIqXxSyiNGmOuwq4synko7YvEkURX9
pgeuRNR/GEiMVThu3USfA437GS86a/BX2Zabh57e0vNEpwG9o3lor5BioNxMVjLHUBfQm0a8GlJK
fJjIM/eOYday/wXd316H8FtcInUobhdkc2jzOJqqATEPhjnasGaIH7PE2oZ1m7usI5AIW8LwMWGU
VusBJdnrkiXdZ8M2hUolhcG33vgi1Ayd8S56qS5ZXZYIpU69L7LGd2onhOUW2j1TyNtYckWX+oNm
Vx5zjtn1NBnNTJCOzQvoGjMIJvQsMEe6QusS9ZiHkAQUYNcrPcKIrvqlA6spW/Bs+xJ+uihOaSmH
fl7nYLXr67hKR1kPKF7vJpMShg4pZD9dpZOPcofx1yh5c63yadSqmJg+xTQXNugbBfoeBUaQDON1
c1zU8PVi1SLRBvTlIJWjdO1jRZa3oOVnuH2IG65ohoFxGyHzu2uaXlyRD0wG69sqYjQjdmjhR1kJ
tdYtz9pzAhUcc8iZ5RAL4gFhOpXLVoTJBbSYPnzXtqn1TVeozDzsTg1ottHancOYXdA32UvZpttS
kQ/5NvuBETJH1fQv8lFPyGxpUEQxtEOoMkOo37t9k9RFme+RYQy1Kt6Ldke2dnsEuPQ2kSgBoFOB
CQXr5qD2RYsKDAVwtmSymxwzYzrHflI++MKfSHELfyaONOFv92+R9UP2hZa4uR5GiGO46XX0e6+5
onKpQ6JUmxx1JbglDPWOjkQyOza9dnbVTivWJ8nUS35/dpfm72JvkZXPFMxBwm9aQzvJpqvloWCi
FvIaB7nnj62meX0R4pyWFtDV3XJ4OGvQVG100EIUDl5hPqzZhiUVx5XnQtFb4iajCHlKPvY4yeKE
SND1s6pFfAeGuRzmKLcnuXdzceR7WlV1/URMfcNcvnByf1uafYrTjIeq4TPwpMpWSs+gWIz9F5ct
CODDUxgUy2ArlxMsPlmr2h6qvomDykU4b1DvAfGZ5LCkCgUcx4dLJVU6Qo9Eem6S2YpIOxjkxEJT
Jab9FjLy9csAbPgQvKWmFzDF8IieqUyjxR1Rs8P9dqlTYCs8fsDohC0QGHmP00zRL3t3JB58QPK6
AAqYPOMXLAYtnayrpFSNmRp8s7f0gsrqavoebOrDlkQWgXBfGmOY1ZIWciL41geYz5tY5YT+rFt3
UrtN5rX03ZFCchCiGb0W5JO87aDHV6U3fgHD7cXqt3kF5g83YPM4Eay9hsJWFI2ko7guWFRRRPSP
9o346kewnziZs9+pP5feXmOIQGx0my07P+sdJH7d8manffD9oI8CTqMia6GzajnTLrACqSthb9Xt
JyGkNT30GFwiAslWdcujrhD5hAD40tZiNU/FX7gdyI7qp0hWjEV2CzX35GbFFPXNwOCKZ/Q5YDyJ
9neh+6HtyRLibX3zew24YPU9F7LgAG/+oEWsqqalMrfhTLFrigwIOu2mPW/btgQYYmYRTV4VFJTS
Wmp0CD6CC0ileo4nJdLz4aWk328k2pzFPY8CzdZpQjuiRBI+FP5gW0PL9JaFeFFTkU82zoJrT+Yb
4/UWuRJwZxgI0mTsnB5v3pZUjYQqsEOd9AzxeSubMymuc+2qZJiEDKIY9m9sIb6DiNPd6kbjK6Xh
gdz4eYQPSUurL5eqVIRSsD0pvIzLTpOVszEPVur5lI/6IfmhG+Y3CBX8DULf2PwZ+tKczxs0d6OY
wVFr2Fvbiehp0c0xSAJgtNM7I+adF+IDKfdyQzQ6+6RekLzeJJOvMLWgo5hWzwWCZz9ticq+0TxM
fSSHeroh7PLmEFORDd0yr+xRcw7Hcj8idtzC8xsUQY9gfsxmHH3m7zx3TpBg/l/K/giI0/n+6gbr
3IWP6Od7JNC/N6y6EbkkIjvEsylmmfXHqpCcxk6XoruwXHAEXhRn+w9n4KD3TDXySbpEjjZn1b5u
zwPPnNzm4rKJahyYg9REripLWuIq0QkFB2LvSoyEIsBrvOFtoz+YDxzgOsi5Ged7QlQlOYZbkrF2
EO9/5ljECdx7Cy44D1Nkf0LrRIT65jlTH6cBQaGOiiMYzKAc7PimE+B0AnNKzDwu42/hwFhus+Fw
L3wnMdcxbIj/Zpjm87cEc9nHv7UUm01HQ31p3BaCv9QanMjCogmv+T4OR0s+ESGtoAirJuEpKy9W
XIq8dXJuzBdMOxmbd9vvsjk5kQXm6DMLHJQpuYQgqnna1Xch2lmmp/4WoKxEUxIPE2yCVW3LkjhQ
xybB2Hc9aX6+xBg8cTW8IruiLDP2i+h3LZwLv0+Y32OND2I1cYJiAFp6YlhpgN4eDKz5Sn62rUXH
eYH8fRyeEKOi2yKGaSxXLMINyJ4/Pa41brNU+ledWX8cH3pFifYlz8eBxH7uLHHtlz1xTTVBRp2R
3kYkj8QMW9JYJ61a9t4Esh6Pfh4c2XyFXpOsRBqaUoP0ThBVC1XX9mJKmIt8KdrK6Fiq27UmKi/m
iAXyyxuAeBNCTaeEf/JYVD6aq1Ne3Gk1R6VpdMorOMhp1iu95dOHBTC+UJF+Jsf830uBa1Pm9jQI
7vZLOMe1XtY1jO7sejSim3jyHKWPnMomQ9t90Ass7StX0PDNuJLWnKDsmCsCvAVRanBvLDwYbNs9
3U4lPtfjrqwgelmGGiMlmb8lOzT7cpzuA1NxPq6hqirhHgX6bpw/S4CEUtApd2xB4voUIF8q9thB
gvCQvDLTOfX2W8hVw7fOsa5Rmek/CIeV8T9SVeCyqUETVYoyrNPJ20rNcyi65puH7GJEdRwJuoiK
6Vf5dKgLJVjf1EBCcbw4ssYWDCgHJx7nlY1YCIcak9VJdZhEuZWkdhiSMJuzP+GS3L4inlNufvLm
4AMah2QE5btvzV0a/08azus8lqoWLVhoWIS/PyNcn20fhOV8XNdeHQNpIrdaSmKmPC1GED6t3ue3
BZ3s2/oTEIXIPxutE0PglS6TlSu88XzOUrVIdtsGnp3ADFKV1DBhSdGND9ILWZQhWg9YiYmURxfn
9nxpFBX7xooMNsJizX7kK48AFwv4xMgrJ9euTp6ROdBlcc4FCb7xqhTzRlf4/28ayM5d6APntksU
bKIjw3bSiXvuMJncAuqqtWWKFv3bUBDllbUa8pupmbKN7nw/hnZskD71vCjrqH0zZSsXoiAOazyV
aY9d0uxg6Wr4Bvu2nLfAfPKQIX4GZ4djN9l1r1Y1s6OXBfMPlVpOGb72tCPXYJtMjLmDCbD64SXL
G7LQOD2Kh7uACJbslkAe/PxskJ3lMZwGZU2CEK1Uk7KKgEEJV1E/llZNXDR5cWNSo4fROwejqWfC
znvlHYfKTx+HiV/WDbNNVx01XnCPD926rs0IUCOc790iv2FWQ+lScQjgL018N584/0qS9XszwAzO
WRExBg99gzAwzAe7krWlBFn+85ozyd/BA0I1SEEXodoeXIi3hy0ii++U8Hs67nP+vtiFibnZg0W0
lHYqXlvZUrNaerXVzEpV3ddjhML8U+SbZajoY+TPOTE3UZFa0ldQd12qPtW7dGhcCxKbcxirPoYv
Jq8rrZVq+V5CQlA6KWgYuf/ydw4b2tTeCyq9HLjRWo6O7gMXxtKzRAyTn2c5OzAYXAWl5AWEG8U0
5NhewL0GBl3wJIat7ZTZQTI5Vvv2aO1pyDx3Vs8XUZOZ9zMPJj8fMstxAwA/oQ4VYH+GpxBwQ3vO
3HK6wBCf5+/t02iNiNAZYtTvb2QZ3hTHrdOcXkQfZixK24JefWr+7a/vf/St2TKaXCuq0PbkzLZW
00oKC1pBOc5CcJ+yBxNGiNXtbPIJEcq9mbZUbvSWWgGpPVdKGzMz7ZJLLjkBrC9yxzf4FdT92R6h
yz9iozzPN82bL7p0vY14rGlm6/hgz5lE08A/eymvjh3NWy39pfa9zU2W0YPq2E3Oxt2jYlTAN7b0
3vJr/ilf/IMhjC25ZOh53PCDSKX2xAskIAms8N2JzVoUqjPaT/ul1hwHMAvO/UbkhNMUyS/iPr0D
ScIj+nMsWS9AntnGHr78rKQ/4SIwqBKuzqa5EuLyuGu4hkry5YRpamb05XN35VVQjwAxYwUZP9DC
ym1ijaLGAVpjCvPR5BzYQSbT86tVz+QJhtjyNJ2PPhnYzGrXVvnyy0sTc3bvjirGclE1nbR7JhO4
W9OMOTWPSFwfQydMrnGWW+hkDbYHYw2/98T9Ezhjb7jndWF1nPntiKgtDmgPOTNFK0w0dnDVX+4I
7AL2RJBYxQLZD1sWNWndbC+wTeKjJe3W0ib7Zcfy9f7LpSVb+2F9RnjYCyPgM71gfBuVkyh/yLZ5
1KB5EvznJm+DoT8Rpxm/V5xEkcPH6dW6tezyaWeqMpi6fQNc7GxZW99ZX0WH24y9KDsaHKfaeaJ/
X0jvrdYqMI3J4i+evQxmZtukkF7tzXFqOXFQSIAiuRTUqsTu85fVmvgil4UFs2xNJf3BVYHdG0fy
Ll+ApJHJVYUnF6f8ofT0SdFy1AOXORICgTMkhRoAuNVTAzPfHEOo4a3FJy0seoVWaNmbECpnOhcP
fVQgP7H84oq8wmEMuNI0b1x3wRENQqxeENecicuU2WBZz3yZ+L6Vct0lrpHor/DLEcsL2w9GW6Ln
ixwQF+cXbJEobwxmxRuoxETGxnm3YZM75kDJ1G4Diqh3LXvEJXmAKDDWhcBczNLehXXV7iPREDK3
NNu1e7a5ijKK2jEVdtWjR2WhUJ+9A/ve/JUztAxFAEAo3c+98iP8e98JyQ39EDuPX1iH2dSDYXZx
0Z4id4ixsr58OROEEWCg6SxBGxa691eBqeVF+uPvkIz0P2K5O9Bl2Hibb4RnnU9CYVtzfeAU5JHM
Z3oss+sfvz0BrlhRQAHXcsYoHdpoZH5rwtXjZGBbjorQwtpRV7/hOXtb/4uZjI/aKWH3ZpsvaqdB
Yi2PwQd0hJHA4CfQTmPECmYire5bxyWDfzsGKjY7O3VHQmrS+wxEP4AigF8huk7XkbXSA0X59oPN
fE8/SHEZhyNP/pBquRNHeZcfrhP4B+7JFmWeJw8G1RXDoBRW+Qlr+bvNB3zaU1hIn9rXpxA3BMU8
8hwOSGlP1t+OHWNue5K7lOs5k2FAoIzhXcRrDceAHgVHyp938rPcCwcX2YOZVgSGJ8FK9+Bwz1js
cXO8VrQIjvlEShxbwbWnCdoKVmfvACLXBA7MN6U4LvotYICSGl2oryo5l6VKxIY5N+2WWIajvhmp
Mj47L8rWmi3uIQSovYN1w0rXmw0KnDIM96WYBFXILuBYtaoTgI2czUGWdH9AkXrCi6fG/xntODng
fQSBiV7COIkqC6JggD4+uKJzwNAUw/VJ75KUoDAd4GmQxTMiQYhzLu731O/cdLA7NrA4L8aUlvGY
zvTxaw8ePwrud1ji3c5XMhANmzpdwGmsZRFx5gs+pxQFTZ+txF+WOxTxl3W3jf295mwRQ2hLrFZe
4vz6/kN0XrTBDt2q537RPPbp6OFywEsGp9YZN0cObrduOW5ik3ySZ4HSUzyjanV48SgoQZpQkMj4
SiwqxTM1th0u7I73o/fnG8v3nikSCZZf0kUKB7JXkCWHUwnZkxi7VxPc8fbffE9DRzkYIPxMRw5Z
Xx+gKBbYucL38gGVVyedjh/r/rwFw1pJggFm8emN74KHLyQtaInVP2kitiWp9vnYJPobl+GDFmck
XM+7GQVW7lEhYyO3CBBRSMXd3740ls8CaCA+al2Ajgid6TPmCKX6re3Wa+oNjPTYXHPAfYNNsy23
ixRawCnAehe11vLM9j+tcq5P2b82SX5S3eQQ6JOVsDx1n/U9dZPQmcSQJbNmccgAUMui+oAezl0h
ZeWUNQUTmAheo24CCmDEahy4hutNqaXYAYYBhNQ2zS8KJwaq/vLXRYj6g5LGeXNgy0Ju7dzPTHDX
vA3PJ0q4FmPLA/YGHs6Md4Zp17CoXWdBn/wU7w6UW3XCj7c3LCTAgReAM1M+/AgBz8mrQvxNw997
uyhk/zgXxXPYMqOs4iYQtar4RTaChePr/93eOiYXjUCgIQrEJfUBYQ0RaghbAkjd8sYRiLIg3qdM
2fl0kuL4RXpWrYmWiBOrJZj2W+9W6PqzxG5tzUjKUdVBjqpcONCHcpBeExSRkqg872gnoM8ZbE9I
QkJW4zhGfMZfkwuTnNQayNqG8TyTOBG/POALxAY0AEdVH+4ykC2Z9qFKcZJ4GEcavIadVNRtAshz
giH/RrEYGumTl8cYq9lMZu+EmlpKyMUIm9/0ugup0OXBE0AE7UoPtWJ4Jl0Yonft2OqD6Sl/7WoI
YKYf27yuJGl8DzrwcGQaaXV8SMLQxM38LZmJFcIW1f175ED28nBdVqvH3qNsrk9Kh/1YCL9uh2h0
p8z4QLO1y6q3Mt/D6yD0NAsdvH+8lV5tM2tS3dqHpyvV3vPtH6Xni8TUbeMgf7eWde4Zdv/z78pP
h0kql9tufPAMH4WXzZ39SPA4Z6M6LgDCc76M70DY1gDzls1EGXvmrofK2bz0THQghiV0MqC0M5w6
gPIsujtnDDmOA/LKhluCutG2LAzYG9zaYi3CA+CJ0B+3XrncocCoHcbBJtrVvKq3PW4DQCKWjV0T
5mWm+0dLFsdqL8qPPPfzxuo+jw9MwnEHO82GOicxinqXbubXlhiV7MpYVvQmjNYZl9JBSTZ72OnI
cMxzSatn41Sz+F+MILKeg7jRz/MDrZxOmyzkXlGLtCb/gzgM0r+BRsd4lncXIhVnpufbuiMUNk+M
JivniHMUWyAg4SvtcFix3+XPUZ+XH1hTcvrsCfHHE/Ba3N4pM23SYauBnvH82WQsOdBybKMZwwRp
IqauUzj/FL3o9p1WTJMwgLhVaWpPmH2vli7WMl+Bwvg/Eblgc+g/LriwnHXdHfbQwqHqbjv8z0Kb
3GEs6aKQQWEJE8Rz57w635yL+zZUIwCurKKbXuPQ45KHneXSECvsSeKuz20UorVMFxf5t6XZI8cm
PeroFwWhDPpEidpm+r7O6dd1WLO5kgw+sP1n+6m5BDXcrq1D9O07unVrBW3GTSweMtckxxPd62HC
xNwclLJqXRL1nQ7Co4W537dQU2BIrM4yy5z0zevH8u3OPs/x06Mnxvhrl7K8xZ0ZJOIH2YObM0FI
cjSgYAhVAOE6sAozc3TYzF1+HlpuHTXGfDYdwyHJexyxjRkJHlyoPrkMkDWxoY61lJLAgn1gUt9C
Lnsq9K0OZQq26TpfzNCs1WQ51sKC32P14/cOq+uqVSAILH6aOknU46aNixKf9nuveWRa/BK9Y9Fd
FVIsKtgTqE8ojdmBYADHDQi4yCMGRmby6wmXZ+Cckjqd3uKFd1Zn0RpPFlyKozyGXFmFpJjDeXjf
03jQ1J+g/FI8w6X/Opb1m1OW1ULcWfAESWVLcfe0hjXKtYUfh8Uaqz8TJhONAwpU4wZ8deH+KHGG
Fp55KqJteqwcdFynT2pQU+f2vLAG7PtP922tz/r0hC9T2RcXXeXcs3Go57ZAudB++e3WpEKC2dk4
gqPjk2PbFzx0Cap8wiAkWlpwvkMFaX3MNgFYaZRGJXrfSelsCfRc5dvy/X7KrQ0d46iX3ueCIIZu
Ih3R0MtX3ke+Q7o2nhfD77ZoXTY+6b6yy/K6t+LndyfKp2Odwzr9uxBCvG3/nH4kKAQJp1Xsfzu6
iOluR+taDaDAuIuga1ZG4Rd31znFx/zmm37ESGfhj+e21IFZmU2yFgpR2eylisdK43GrxxEyWrZG
92XIbHG4xcJb6CMH2tsdOIZj/AULQzdCIgFLcgs9ulzdWO9wIPpUrQsHB0Te3Rikhur1Xi/FaE6i
TJrKSOjBREreZZ9vpDEk2702EMJ3u013n8n6v/R4vpnmvOzzYepeKQYxPeU6sTkzmrUPcMJACIf0
YlMQdHuJsAGVxAMTSBd2WvmpeYJW11gDcLiOTA0T2bqiEYS+havGqiIJejWDXlC1+zAivA8ZSPPO
HiMkg3W1hTHPdDqHgXyeqlw3sVFIcDuLTBc7oOwBR0LLc+TP2PNFbRtQ/og+SZdneRm6ZaU5W9II
rTZCRerXRakIwJGoNt/kmr1j+ggFvucqm+/XOFrKu9rjhGii1ni85DnmMu43Q9UHN8hmRcL2NzaZ
5nfvsttntsF6hAplwBjAaIEOFEkv7K1PaqjIAKaFnQpViRr1beRenvS9LdJqpdGqwQp8R0cKtta8
GjiBFDVKxl1dUHbh7YrZOVnqkF7q8V9hrWVd6SmFQ6VLS2YJlYifw64Oe0fK0vjbLkjVIUCz1ZgO
onYUCoRwu7Im1z0Ww6AZrLPVex1P09hlmBdHjP/n6KuYuOfqeiCmnNI16F7ARC8YY6utrDZ+kjWV
PGzvMGlGYTvOKpuB9ms2ZLMBGhZEVNeQQ70zW7Fat1Oli/VbGZpAscmyPWsqRntHrFV0LgJX9UAt
C7XDypBEZfiCiG+nMb3zKkS/UOSrEwVz0TivqgSVWcCqLRoMDOatocukNWK2NLVzmXZcixQnawMe
nsugJQ0iXy/wg0sNBN5yk44XWPBI1itCwI6y7ueJqasxlhpozhcz7TdJWtjB2ZWwygNjBXy0XPGs
eay2WhHil3mHG53kYUA2vDTw/cp1VNtR/Oui/e+BNLKv79QJwBtDpAbCBZ8rzFrVOEa9hfyTufNR
rIId0Pgz+KYeXTkagWS1RDlokC/bth/ryRJFY9uxYimI7qAzwnNpRQxmChI1fyn17/GajwsAn8zg
s4+bb7pxOaa4FZmbYyL5LK5a8WUY0Kcu/pCZ16uXq2cWoCFJVQiZaChiENhXX2grWOEAtlpAyFXQ
TzJ82/YPF4jy5u8AXoVfY3mOIfpywJKOgJmpkEjPUxR6nJN692/j6HVZh7HCKTO3dM2tGZLx4p3I
boWbFPaMR9lKlpWb0ajB8m6olHRvi2JkYx/nhL5E2QT4hnKb8wzF5u63a6RPGPJPTb8GtvkhM3Gn
O4IUp7dse4PahwM3VQ+0nETojnHck8+m3+CHb18Sk1fi3nfbF3o6ebPc0Vzp0NIUqytfpWDZQJew
eoe06awxQDjVuzyuqLpQj87XPmiDyAWFauYD6+YMT/yvLOt50UpDd35Zaz26y/14oPf0Wn34/zd+
FfNuL16fgITIPT5x3v6UgtnlgiKeGoUPBEyRP3eXqd9teQU5znrCSjTX9tyIFR52MjqNdPBv6dG1
4/+iwJZWy5OzlYZaV7vl0VBC5Dsh1QsUG5k1CRL2MP+VH45XKCwrG4JLDDwpAul11n1E47cz+EL8
i4/pByJUlgPkW82KBpZLIY0Lvb1QeyPG1ZttHT5BHu+pFacvBm+8SmK0PxJ+7UT9fXxiFzReK5Eb
bhvvCGuYVFBLzW18zkr3DNrm52YfZw6nTclX8FjzLE0SNQpbln97lE/794QJujzhNjkRC+iOXwMA
259HiwokLyoEZ1ZKD9zFm/FRLaa9WcV0NFDC51/y6jeN636kDWUbfkQ+M7D9UH9VnA4/YS70FSxM
dr8ISOma11Z5Cb44JcHH34Gw3Plm40sWJiNW86XZZOA1f02iz52kRRRnlZVD1OPVz+orJaP1RKFO
g1SdkaBNsfgC3oKUl79/NRbI1a4VgM9YXuhnzw3PN46F3wrcsK+L1L3C7yYEhloYRxGfqCiojnqN
Luwd22V97FCloXudh+TGPwaVKD2CfLTeeLOWt8jzmOHiDpj1Tjhh3oiTFifmQLCl2uw+6+OVUOWr
UdsYDJNtRVuiY7ivVsAzApB+wtjDXtIZCluIvpz1pSTbjiqx0wJiQzOlNuY/23XVham8W5yrPB5F
Rrl9h4k0PtH36yzmoNnryp5ycQ+rPhenjDcPW8iY6Jm2NJf7r1ImO5vVs0C7Wnz+KNqUCdxykh+c
V9ArprKdQBtGS7nEhKPR1xlAA1briZjY5Tmst/6e1GVC6lGgvk4qC5mD9Zu1uk51m4EUkU1vdte3
q3MZPaZOOrDwRnK/feuTGaaXfsCIBKbmJfThrWdlDBK2CYn5C7BnyfDST2+wo1ansJ3R3itMzzg5
/AItMmmlg926+vpkEL7d/NDaLXbgyGwKmGjgOAFllb7IUXLv/eqcRb+w6fzHoEmwkkF1qCCCIbMX
kOtonq6KmuLwd334T14ppFBYNP7u+nOVyscUc0B8vBFhuwq3SgF4X80tRHdmqnmMFJpAvnSAE9Gt
3q+PjeYiWBF65q7HzH66AA5KH44cn3aQkhjayMzvdsbvPhJYLBlovXr+uiQIZCs43miWmblsY6ry
CiIrP/QrhgEm5iW1zTHJ5XdlwG3eQciGmhfCJ1+W00loJFxWQGcHAlJpBUV34JIsb0QW0kZtKKMr
vNPxY+2g7mnHSqAInRsqGdGnsPYZ/ZKo28tjhFG/EOQMHmBFI2jWbprs4YRIX5jm7GbMW+Ow6o62
89XECt4iG5rDHtiyycD0w/f4M0grrVpeDC+sp3nMNDsMas1La2bdwd9y+sNNX3KD7hXrdlsXy+4I
7I0D4G29WwcfzmPP9hYJbIjvBQsQL0OMRHwzLc4GenZCGtxdosgq3i7lKjN5mHKIWN2lqU/b+RNC
/6dKIJkXViA22sYYI7q7iHaOvHCbEQjqyjbUhWPwYhPlf5+YiBvI4pNLmTiQ8faiTeBhbsTAqFYp
PpuDPvDnSnTPmE69kxn7fSnABTDpsA58NgrASXRTPteN6U/vXv5OCuJNIc+IH++0GMyqR+vI1KJe
+hkl9xG8/3Nm6hm9kAAM63OFybG/BT3ROz+6zTV0Qou3a1EDnYz3HRGcjnsooLE/c3nao+vCqCjK
zIMJoluOmQ+tNQBKcarhMhZQ9NmfHHAfggoQbXi/ZgSaYGfBpK4AWtwM95b77IefFljyLXVyXDy0
fctTF8E0mVGkujuWYJzGGSeZWMYTTs0taVH5m83aAKdF+uFkq/fvQUWwZUWeyYaIP303RMhIAa1E
lzt74r/IIijJ0zaIXnflb123GiQdygEJqn+ZYAYir2Hs2yI0+T5SpspXhQu0fXhT1yrhmNo/jhTV
ysj23EpnOAORbnEeZI5bKppU+R6UksC5UfYKku4q7kAMVia/BlhnDVhANn0QaCNjmyNKvqbYblR7
CQcV8I+Sv69yPfwKSVR3cjApxWUNi6ukOns4pDKV3O7ZMtxqin+ywhRTBrp7kcdkInjYYll8Y6KD
yCI3iUCmupCPOmJLfDpE+rInebmDH8qKICgFhcBDiUzJkC1rRzl5pxsTzqKyvYyhfQ03LOS9wCQ4
72pUvIuXxuhV2Y/yNqCwrlmZ2mh5yUKTbzx9Xe92qGuFa3hkqWXO+mgfoAY7VdrNW0niUSk8qF74
7aEVL7aEXu3Tw44eq3dyEKwmTZYgconGiEQR0RbWODjxVk21qVmby1pPH87cuqZ9ESwjGdVq0njB
DXBktc1sAwahnZ5hwFanR/pYSlhvgjX/u3U0wyY/SLSE9Da2GSR+LUA/r0aFjcsXtI82EGm6zcKQ
Vxlcj4VWloZm62B7QnlNYUHh52S4MaB4nbkd8T35X0qwXfK040s/jOEmRSnzMIBCb16Ajf8V+cKe
miqXD99PBU0u6b4/FoWKq8KMe+0Xavm1Y/zfogfy4D50x/BXYgENYi4MBKYtgiygqsIoS9+MNLcs
sYgoYcavSizIQ4WSmoeaTvq1jq6HlIGlpJ92Swy9YopSZBmU+28eoTDfq0cyOi+ns9Kwj6TUWzHd
wYdGoW6t4aKetRxqU615RkWHmY8o+b2imGbKlW+TqyT+4gJzvnotSokNJSH7KPo8D6BM48aJGbJA
sbuX1X3FR+f5NykcdtgJzjDez94kKJknAOQGLeAKtyBns5ncknHiZpGVrOvsxAkeCLf82P7SqlbO
BtVl81hozRTp2EKVsiSL6Emtl0IBkWZrfV9pCd5LSXcKz32QtL7vs2g0RllS9DvlVogLsVkBHyBV
Wrjff+KkXAHbnXE0oL/b+13yGb23Mm6gR94shrB9h0r3MB97zJLgdzstiWDfYe1DzxKxuT0hL9Ph
4ewiBTqCMHNnvXAcMNVPqAia4II+QyBtbgjWWiZUvEG8W16oyiheIbysFNXn51b5JjduOgr0ZC5M
jjmVAY/VWgG2J9rVqVbcFiXZB0CVub4P5H871Da1o5BdBRKJANFAbINrwwtFkTAhctUCbfrmQuOa
d+04le+4jcTtEMTHVpVAyyxIvITI9kSrw1VcTEBDCrc+MUD2tf3ywS2Lm/Y0ekOE5G2JvzEu1x9i
p3fsO9Olg6sdCq1uQdcsquzU5+QUKPn08UpStbwtE0w95V23gVB9kFqzdkfIvCBq4qNmD4rTEo9i
w2WePqDfh58iz3rBXirsXLJLnrrs5VDkWzVVGQ2j2lDmyIfVDYQMRZJ67NSKkhITj4Gu3FHzmy0P
VmaYnR7VS7TtRUcrQkEDsSWA9NPB6N8/Ewnj7d653L+7WQYgsN9XDMIa1zy5RqE2U/Z5bCzg1Gce
1gv0QtRiPI56qy7Hf0Lfix/soU/KH6W0aIC0qAngOSajSHv8/PzUSgGSMWYy21zruG7Mzlvt4Pd4
t+ly7HrgrtelYpmX03f/e4fxcshPcWzPalSxemGvABRhPskTxDj5mciOPFukiiL8uezW96WAo62u
3bYcPMhPfVSComkEaNS1eax0CTodBMGUGOR6u75KQGYXeTHzgg/wMy7dlVRBArTAlgDEv6JVHlme
VVG2ZmlFsXFFKx/1vSjvNSC3P2q82WAmtyy0cA7pWe3UwRia/IUcXsiyrj9glkrtvIf72rhaaMhD
K5uqeW6Q/EvhYOv0VjPX6prrjI+ZYRBJ+5R8hcTztj6OySJvYuJqrgoWQtm4VPQo32sXat9iZhtN
tYHP6ChMeisrFrZ3vq9HO/U1eb2D/IFoAb3QYqN/QrzC2iRO7LFBCK/r7OAz1Xzw2ocQoPtP4eOi
cZ8UZi6mlJ9V2fbmnZEGCb5T7IpGxQOvFwpazsOsqAotl1Q399YjlrTVVPCG3DHkwZvTWjWIWwGF
7vIx6o4nBpdT0861D73pljBDrMMHxBgD177t5d4btKRFiXSwQf3CqyM/SHL9tl3GlkcHbwsY4wOD
6lz6k/Z7Zdrx5FqDCUdAJtaeSVs6VmbmywPnAGantpn+ndP69Lp+qoH3rqgzpdXYiizB0NMQDlWL
6abJZZ8ANgYPEqTdLOb/OC/vTgP2NMRrv+cTNALphaQuAsAbg7WpdjVlNLffJ31RvuDjRixreSPA
lFbquf/k5o1CElBZMJE53IFhHvai+LldQOFFgYGHj/J7eoEkSGQryI3hXGS7zJ5hXhDbIVVYJCWr
Myrme4aWIc/iXWy3qkPVhiOthLB4Ounhcfd/6Lr4Pg2HzkrW0L5lrpSw+LnnxTPeTuZSzNqRFyc6
s8gEwvVvd3vNgjUQ+IsUfS33QnXUASsCSXJ85nxv12zzMSMKzmlbFYwEnQ0h+T5U+zm0srmr0E/R
i4S7RGLqajxxh2lc2PHR4rWaKe1a/L0uSp9z2UvJFNjVq3CMu2L/jtJ8MbqnV+RjP6VoBw987Lwt
JRiniSkPnaDgoFwbOo7N4/khgK48dpWPMYN7/GIrTXQdFoZuReYw8cEemOQ0dnGnO3Wbcs7VWDa5
18fDp/s1JMHZXwMnDQEAkyZfXun/SZGs3AbL0qUA7CNPSr34aQpRZZyJCk21F2oshnM6MHky4GfB
VEfimc1JdOnYeRqH4sNjb6tPecbnb0+bPbruOGbcr3QhAWj91k4l616aViV3rv7CpkZ1QDaKT8Qv
ffR5XYJY0Eotx90Q6hYDj/+hJP6cH6dYi14oc2dnbK/0L6spkZlaOOqwhpUnxzfVXKsh+GxEFOif
XxI87CxNy88KCyuNTUKp5/MxE8N1nF+rLcS50A58SQnvjeqtv2PigpbN+pisdcqpWewx8BamksX9
9cZAu+esHVKj/TWfSBcqdVodcVDruHwW+ubcJdwhQOc/8rW/oE8VvTDVNVen9X9QCybKx24x9m7U
kgxTf+KEhKUjqv046vQCqnALRTBL2178SMllDHyPcM0ZglOg5hP6uA7ooyviep/rrrrKppLQFQM4
AQ+h9QMQPjMic7o5b/oQp53L9T/8YgCAuuDsnQfe5Go063MgUZhZ208/ddn0E1npL/q4EGMf71Dv
BUdgHNLzJOX1xwI3hEG93NbSEkbV2h/TAl3pCAGfndSpZo4iNheM65STf3muBtAj0XXarEWzZpFG
xAocVTWToHJmFwEKANRmOA7HNtUzHhH6hblBzAbwGlKaOAoclRxutCf0YIMWnkPGLxwX1eNLNPt9
WZ9ConEIZLPgiKwUyymYvmqqJhXhwcwZAnXHwhJ4LIGOo0JBdtmUYlQjJ9l6W0QS0UwhvmfQfWRg
hi5hfvV1y4iFGp5iwmB16Lkp9cXIJP/WNXoMpwFNG1GcHYPogzEfCd5ZvOgYypIVupBIGlIVWvP7
TRy5KuRgQsI/qgTBKZYcH+pfQAGdRQCScWGTaowJ04ReNTVoEdSeGr4QofItUWaVXaEEDoKMRxoR
mePDll9YqAottP2oOfz5MGj1WSBaQ64H1w4VHg5BQR/wTFmgMUS+5MQ7AowBPg+wXNP9+BPgjGfu
MzhBrfaoAG5Hrzb6Si9PwdmxKrXE2o/fh1A3Rpe6QHQpabZG/85w7utNlOIjkXBv1w3W9DYLSAO7
zUDynyXnLRgFt6AVLlViR5+OjNatyhDKwVqyOX4rSmpHBkoDKdtEXOcTa+ZkLDpPb458ZZpJbg4y
5liL7pIcaQ+c14Jav3VndIEQ+zXVdF9BX9qaeNhN3nzecl3Ghy4S4Lvb9uLGlrMnXkisP5eQLGLe
bAciUTgQQ/DvKV6mERplCPSwB1jArhXRxJoJGTg8iqoyGbClUW9VaIwYah9vr7Sqd6bXch90VltB
8CvPWdS9nqjs/IgbrjKXmJzu7i+cBLkiGnn2P1KnEQZgdWDK2JTOujlRIsI+h2jSzBn3E7XP3b5E
0Q0POLgc0jxubwSYs7w281BWSVw7dsn3xAjRKHvixwLwk4eE0122f2UGqkrz6UD8Cok65rka2GTy
GOOiYugu2xe0cqGZG/WJ96MQEfGu6hP76HHZLjpfkPb4jItnCueycZNZI3Uesiyi2n2AcMW2vaHz
srwEBb3HIodOIf2Np9KlkVK4lgWchgJa1gKQ6LXUOJGncd2cOWQyV+stTCbeTWx2Jlgy6xDrNv7j
naORFEq23IL5KOoQP/TpWtRWBCg7Hr5XQ5a8VHaf7wEQW4U4p27tTFpdmaZ5RshkqSOuE6M/HbJ/
C36bShXhPb2xx5nqlH424ECJAQpsufqcCJxqqpg4x7e+EceTT99HjQtD+Dza1mTaRI6NMsc1DS/M
V1MX/tFiCQgeOvqWDynF9SN7zlzFvcNLHXMyKjZ4Vlyz30lMIYDvK47Hdzk5GLv2OAidfT/mvP7R
4mOIlQ0T5f3M0BPUXLvElILsM6h6pjYd/1ZiHJ8qcvg5yjirVZ/TVA5YxZ2amwLn4i8f8y7XrNwi
KrdzGLohE7spjCCapuGjAlV59P/iDLsFydKqGmv+qWUL2ZMZVoh9zEuhuwIorHGp0vx5uYmSnUzl
K8eE0FzAH2SjQYAOifdazvyoHap7E7fzkOw4E7wGw57g9VPSc7UHFFQ+0uPtgw65ncFDXDAddMpZ
HT942Tq7Vr8JXUwv/tvbpkBl7Q+HSoe1SuvAVeR4NNYGwC+o4ju+xHCy9CalaHkzkXLAx+4zBqjV
gYQ0MaVGZLtBL9IyzWVxPipcP4pj6pLIUERyEv5nZup1KMn8O1MLNUYobcQekQaXM+TvSnP1YS0z
3nUDvgTG8mwCREdjMIOQAC1YANC5lWIDypXWy6JXfRFd3Kem7ihwemzVA3GoA5inOrCY6qOpI6Bs
7QLIttr15i0BlWtJGoBuC6ZVy+ID4gbrjYPL9QYBtbLnLeZ5yc2agonCinU48Sww/bK1rFX2DxjA
3/yHLxnER8fn/UVS6VM0gsZI2B/fZfbfSAazrD+EHGBxf7hnFU512cBNA+cjb1zDDbL8i8iNjZ0H
VGVhDONR5KO22jJA2RY2kLLmwpmNAMQ7/wxzCMzQFf73jbarY5Hi1QNx8b5+hroA4T9tLzG5u3et
FRF4DisvA3qSqs2vawxtbTOJREohvPihF/RSDseuio/xMZrpKLv12iYIHMgr2KO6ye45qWmgGtJA
Yawq24JtmI5AX/YqxXwIGZBKihZbx8CYe6FHeO8vjcuAFSXoG8Hvi+XAbKnBm+fWE3vkfjfx0jHW
p6BnXF7FdBez6jBiHRdFQIy4pfBs1Ju881JfOr23AqiuvGOa+aZNM73eXnGK/+GfEQo+Z0yVL5AF
q1iXaaAiEdIZe55lSdbWgmW2CIIyOQt4ZWvOj2H1s7shguUCPaI82vkGrmYeSc9VvDIcSaK7QGCz
ddYqoS2+D0ZFO6W3okMHDJCyCMh0XONgcEM2WPVu80YluG/Biyi7Lh4MpKDwYorvIi6kt6loEl+A
PptlBMy3IhD7JvEs0mMk9r8mAeP7B0B2qT/NbTdP/79q89GdM0i6ngnpVJrfd/vaTE/5J0bi0T+0
RgBweAFg3GLyMNGagd+Q0Xt9+wPmyEya/UUsysngeySuexW3mpOlY47q4FmXtrj6PQCX6QN3GYiC
wO0FAo3tOcgzo6YOhJA7afhelXlP18moveWm7a/yLDid9MQf3Mnjo49Ly2qCm8MiBqsqTaD63qBj
meigrPeS1HPG21ReqqTJh/QprQnImIyRDCJjmICU/E8N/Qy7+YmYgSoMkYsGH1PEnbVSHBo04yuo
jn6X/z/oYNFlCxcpdakPdSBj+whcyBHYUK6gsJj5jqAF14ZBBzNvthLusuwymQ+N4cchijlK/d5v
T4Ejgy6fNkIHDpraK4Ge37yeF49lvAxqWaASorJS9A2JgtgGJf+rKRr0hMsjqXADB8yNGaGuX3je
c/GR1w8eATjyZSFHwtBp9bvWL6X9G6E2ni0sbFo+yTqJEUu3ga1h+fbfm2VMV9akvZ2IorYjmJOA
f97rn501q04v6LeZkG03X1Vwj2yQD88rngGQa/Misk3nSQgstZ7meht5ZdZoithMwtYk8xkPwNao
hLLAhq+Mp0QydrFGK3pogGLpKTiTsxoj9bKWWC/tdP39/+sGzY0VjWZpNVF59fxpsvunaLnc0/6a
I0Smg6SmN1auWzxh9Jo9rewV9q2fJ7c5IkKfdRTKrhp4CpaoISmN10D3pTnIuVijgFcL4ER8UF+/
ynnBISCBYLXm0SlFX0UGqOxd3YXHZvgp8WQiB5VS9SLVTksSrX/8LQCFQgloKCUVIoGPVf2krZRB
0Q25D1tY05YFLGrrNocmTD2RK+3aRE7pRqVjKcqzFdFwwOmHADdJv8lHnFk5f4eTE2RbAEOmkZ5A
OcZ/ahCW8X7wn3RzJAHVKvuIGHYzbZ3gUNjRiFHj9CGOBY9nFAu+RMtNLAlV9oRKsrxKZbs44pU8
EWKnmBpiRfsp1vMlv7yIapcXa8mMloeIg1hErmDeHZ8MtIs9N4tNUr4gipTjUgTx5YYXPctXGVPl
5qoWbnxv8rmS7YlJuvbnRhjhlI++YG7rkiWxnUa8WAIlVjfFNIZAQ3d3zW+lhUHjm/rvbDdl78u9
qydrAHreSgv8d71RJIoxbuqnLwIFLM/mMR9nMQyx1f0YEYwWzSu1+1hKJWZe3f4HsFHhqo9ajOV2
LgLWiHvXz/KZA9fVEFjKuIDTaA6bRQlfKAIuBzWbXalwQh56tVJTNoCYNGFEd6fqMJjckmhofbtq
XPag8UKyF9sGZekN2mK8gxWhwRkK+nnEWGHRrs3nXXFSjrZcQ/DUx7ukg1Nxu2BzQ+10tPO5API5
4r4Foj47yTl4poE7a6hGUhYG6pp8M7+PzvEUj8aqFjBLhwXg6M0nl/xqKaVcHcIXACps1sMZb946
oXn7Npenir3bFuKRfgMYxMscINMVZF5Oeqf14s33wqW2+WebULVIaFX23yXsniTuDvOZ8oM0j8dl
pxzIXvjjWalR2WAN1Eq86C1itWtYOp58zKTbjQWyCs6fBS5fuQM0kTKkhaaISNpJUghBFJIULLac
pq3IFOU+OXP6+ZM4Xylp6mGLIl2NPLGTZC3Fxvp7qfH5Z9czYr6hGcOJwLFDCD8jyf5jC81X35Cd
4TJI1OvOwSvoPlGl6mfUG3zRBKBmjtnpWPhj0E8y9o8POodvQ+WlTqhitJXehZTXaHjfIHY3uZj+
Oaw2DC7oPs2j0nNZErNm7NWgZ7lfVqrY9jlGrBRerYhkypGZFrqQHj6RaHfsfD+TCXFAKskkFDTa
KhOVVjiPvkgf2eNiJo3KbYjo9NzQbY3k+TY0CJD4lqlMjNsEJiSOZXFrWqD0Y90yahHWsdNZNLsr
WuwyXctqH+QQRagZtwCUjRZyj9CNHHki2GYL482bpCY4YyGi8Hh5Wav4xZBWYVUHpT+eNrqhwy59
EHV01gNYgYWbKm/eeT1lck4qasAzRsyHQpgDVOPlbbnRMBkDAq1vqJf4oS1vbcfrcRP5TTwLtfMp
MsiCRCueuFup+MFGsXp1Mrn/NtwDokh7ysl9p/FBXeK+/GyjLbX/1XVHap2c/oi5fJQPct81Ux3n
QHkHxNm4Kef+g2nKTa/f5Mvd8dm6dViIL9lflGmTw5vWpuC3Ermy3AofFQOnpBsMJhHyU2BAtmIo
e+Z3GZdSiBbCml1+lBFq3uzQ+N7RElEaAPjLPKH39tiXgCdvOIK3TN/XNabfrSOLV+o2JRrx2ro3
DIIeIFChTQIh63FbEcM1Pvk4YcUP46G3QnoZb0dzFPv1rSCx8M5b58H1IatoVlSjF8aY0kX9esLD
LrElwPnMrBsP+TRwA3l8PgUQ7q/uSDu0xAl1Eqy3GiotVbrbt4J1srgK5yMlUcSaVSIWiEi0gVG+
cBZNGhl01YG47R25GGTB0B5rKM90r6TTpyj36TVoIGagwgiFyjzmGmA4zB+c+ns9fvUiJY4ONKpj
XBZJF22Jn+mjORB5wKs3I1WFGj93/2FCjPMsb6kmhinsMH/NktAAuFOUT8//rmnIFFLHlTrIaSsP
dnI7zegxaQ8ENbwegkyDdqbdKg6VbGZ5zLl0gY4E484jstYq4lAr4P6Viw3fgaCNKpiybEEs9Rtv
3cEQtA6rNRTwiW3iCiYpjaEKni2O2G68s5fH9s46pmYrOSuxDomiLjuDwJuDx/qyx+eALppjpvmn
xOJYv5jRI1d/8L0Oqw1HZRoG/6ZH34ZWVECmIWROeCcyLpqWlBFAJlA/0E6yEv9THb52Fv3Vg3x+
xNPo0AvB7WaL9lMCAoOa2RL5/uzgfQsMiqyj+97wMIyCfH/fDnugqSEKY+fKHlvKTO3NUfw38WyS
OuN4ut5/9E90hmA84nUe2tRyPIh96i+yA0qQvJ/Y1hr/RuMUGMRFZNszITVPFQsHxhgo/6BL/RXf
MUWTEQDV6Xhk7IvUyBtVXrXUcMmC/frbAoFWpzZ7v8fQc5hFyqlmh8DZgJ7B1PBFkpLsZ6nBxzow
OTym7p5oijNsBJM78XG7BLyY4mflFoBKRVuHgAab3ZHMa6yrgIcVrWFP3BFGExQb7Equ8d0Ksdlp
fI61Nqa2zel0RcuLzEfwu+yMkE11kuKK5zkB6NeLwwdIKdw6F+rv2jBdTPreEeGT+EJn7L0kUdz3
RnTsW1q0USDQJuyDdiNstviSBIYIKMZtIVmlt67AXkvCH3V2MksPjoheme4HjHnlqrnq6RTdIED6
8JQwxZXkAdXrhDTAncunKNA3O9xGqAFI+mTPLX5h9kqB9hM+9NmMTMn8Xi+92BRrIfTLjA7YbWi7
QxnQTZkVvA7+f4sw3BP/pet1cQ3kg9JBUrprXqO1Ltr9iQ4LW8pXHcD8MqFSnMNQwxddvoB5GYr1
n9tyB9XkmViajLopNLSpEtNDwp08oYgHxUMyIF2mriXIW97I+eVhj+UKC+DZi3FQwUWQrsvfLeEa
CttH6+2QaFk8dJ+MZLKzJCxx5oPMiQ0L9f/gatddp8UrvDsA8xJXfCRu6kMzhZsSLhYa/fYgjv9E
XhH/EfY2f9EzGvc7MdDAY75fJgN83ZdGMobqJSIKmmMh/MFt5RfZOOT/IbtZR6/hxN8gu+g6iVzq
kRv7Tl+Nx97wI76pjaUK1NCgD58ocm7FfrbYYWgMugrYQoeZgdBOZlyH6c+U51ATVt1qRF3zBk5h
DkQpBezPU0s1dU8uo76ucaVSQMOdMg9LAnC2fCUATwNc7eOmQoGCAjnWuWPavVgLsiH4pVMQKntO
L1uvdy91dzxxsbjDBbvs01PBTRuVfJk1MB86hFMO6nQD/W8DslsFP64dN6S9bK1ceFNnoScvuJYj
OR1/+GttHwHqEYFn8C/e1+xHyw8XTte62GMFXK9qgjnhnJx5uijoO0aMlvgy6jURYIVnIMw/7wk+
SEfUQ5N3cQyypHyazWRah96yV8Cky7rAqEThi2pypGMSK5z0ZBQ3edHVG2V3F7HJiMz2fV9/HvTe
e4aRaF+MF10G98L+M9X3qfwx+5lUiJ7WcvXSHgnMvR85+OaZB5UcEQVvGlCwIuMdmmdqIdnekNfx
rdApQw+2tOY/C1lQmrT9ozBkz6Yxu9Kf2P8b2AbGEsGcD8ySDVp/QEP1CKYHJ0IOz+XWtvMgzcyD
p7xC4IlwcEhTLL6R4VJHK3NbldulN4W2UDUiAMCHIN0dqwy6YZpcX9v5rW3vxnOLFFPr7NsYLnqb
EJbpktGleMcBd4OELrd5vhP4hPSUA2V6O8ZtFrJ2WrIjZe8skrLSL8abmL5/fV8zdeh20g5+ednM
LsuLw1LhvLDEvl/td7gH8vRSbuJo/DRehZBTb2QVYzbeiHKzTFGujciwrDM7DXgxAVl9ja+oqq/J
ROvKn8HzTgWV9nSZnCaJUkEh08lK6/ctwr+KzTSSy877eVztl/0OLQUJLDhZZjys62vC4O2tlYt+
LN4KNfx1tUX5SentKHlZwLpUuUkSSlG8pB7BYJGstK+6CdZD6hBqaSZJhgcJ0gDOp0b95RCtJLFJ
QmSHNuQswG6aPTA4EH+LkuwUoZ2YImgqzSHpGvhxj7SlEbxpYv6F9O6dRbw4Ro/nK6/M55hNU5Wo
eXm2Xx4RP7kFmFzf0gfjggxWp7/v0Iuyzuu06e9ONzKWszVB+/Bd6Er4zc1GrG1LhlisRHlEBRwQ
awOEWjDsFUE77+P41929+wcqmRxe5DiFZQCKXBxOQCpsqiUSJwhpmrosEBbkX0plYIZiSfWaDMkr
jS8vcdr9XODQvuavCQnIuIDPVdUsnWX6qhkQgEyzI8YyVsSnEUStKouz9j6z71U8PUxiVWWEzqeA
WuoXqVrYaLsUYHx+qchzurKXgW71y04NUbFT9tXxeW06LxZbG6Eh7lCJ5vDENwRLmzpBrsPAEWfn
0mY+ptExEJRENioNd7nn4ggC83ZOfbUWRZs4KgoBKGI4PDxpErzKqiVJAkJQtbaPZn7ZifEv46lJ
pyJHrSgV/BJw96eUJNTP3m3G1oP70o3120ddpnIkXdJJPFHHW9tnWL167y3pxnQreevRxAhrtSy4
XJfCVdsViUevV+hAfczscec2ZboUjYHqxIWj5dPfMNkFzJnQA9p04NXSEpDGOi043MY4F8aCGaZk
KWqtDt2Ta5LgFcTuH+4mjlKbYTo+pkzeyx15cT5HwIGlQxKGGr7g2pfxCL4AxFZOGt7TNixy2Xyt
OitL8rDKjj/35IyjJcpO7tdOCxAP9UTmKgQNrOTqnD2vMIyNfrzjwrKPA6t/haNv/us99OBrMXvJ
4msR4guT85/YUeqA5S6YaMYaY4qqVukVPpUMpqYeNPLyAllSrpNA5usrPgvt4Yh2prF+tlNZbDFz
GC7Rp7yjV8YMIQDUlBOM+p6tMo+c00RyTHoQhX+qvtCM5w4+cS6dj85xUaXiHaW5sks4V7IbLWaG
joL4F5vdXFXYQs6meZqwwHiN8O7lacwhiCeg0T1R4D9DTIGcPLVFzSVSQKJfhuR51p3Q0R7+3xTg
p64JRn5L595K0eQKYeyWvvj1M1KWipxrHUu8ZA12Vj74o15CC3jD0+NdVECtLnCwI8hdgS8SQkeU
vRWjEVo6W3CXHcQyXQZcIM7An77so2OVo8UQuHlVCOG4nDRGPqlinHs0YUvp4AMqRLRlqpXwDj05
io5MmCLYGGZqCJq+D4L/Pp7UodoCwfkps4W8iGDQwjjUBeVvoNBJp6KU0tsuvLahElSVSQca8SK/
mj5V+oBvHoca3PeVAtuPx2egvDJ3YMM/ispN/DWmgTjDCaKtDoZMz5W/HShZ1uReajFUcE1BokTx
eVCLeO+nMqSTgI8WSFN0+jC7SJvQtRii/kuA9oZ4P402S4uIiPV83BbZzcKU3SHC3TWc8exGAQSJ
gP+8ifDKfxyFxDt656ecOA96H5teFKBShGM2+IIf+s+2nqE8kJhswiyo49aeGKrYLQEnmnFApaQa
N9DRrFrsEVjZwUhkhaEFUEr/w5X2Jr94ZbvzN2znh6Pbu4jMmQxa0Er2Mj+Zmz8clLc5AMuZJLhq
xZmVLCQxYm7Pfh5njXQPyq0DzpPOhkTkF0USNOWv3Nc2WGOWw10nuJbvLsqvGDmvdVQJjdhLWSxo
y75xvUF/5286drpl10ZJU1FjTMHnSIrs3KC1VBSyDhYcq6M5Z1oR3SKpfjv5pjbUhahiCAZG1f8r
cU8sd6qwMMD0f7b2vDpZgN+lPidQid1AvGwcx6coBmEoxsDcaO9kV1ykQTf+0QkNbC+HIBWSLOWz
LfnMmsZr/ehOBJevykWucEZtVgi2ixosUBzDHX1GLGqCJ/uMAtYh/nBY7OBxY+7A3qUPgXgtvBll
pej1IqurHShcZ5g/8fGgHqfsbk8K/8/c1YzSZaIwyGK6W8nvG2EfvuaPgr4eD0RsbE7teOO3j6ss
rC5J+DP2jcPLLwQT9uyZD9CjXpvDFXoyh270yR8qw7xSMrf0ILkv4wyEK3PJjVCZ1jN8INWeeADY
wSNsZwPHmE1xWgJjD3CyrktQT3a6Xs9Kutch7Hoekpxm4TUhHRuNQ7iock+TMz2vhvoa4RdrpJCQ
u/Ik2QcRqN3B6JImgQIVZg7cJWZZ34gSFBgwPSNS6aEeaAP213e76Jz2oHIKtaqIJHgC1mlzSqTS
FIRdQQSwTffgrIFACLyh/WhlfvpJhDOCgbhvXXBqDlSM534kbPt0r0sBNEOWDgLxXl3NU6U0ESdD
PCLdM93JLokXpb6AjQ/8NcPhXId9zZznqJg7H+7dEKBUAinmQwEdUKYOs2taaI4UJtTubmVOYRAo
x5iaWOkMZuvpjfnqbI0YP/xChsLZkz9oUGLyy2DitQmavZNd0fOVWTmwWv6dEknlJWoo8IPkDwP+
hT5IdTmO401b8lC2rCWBHV5MtladIVQ2ZZNWf6ndoNE/o7fQ7JCUHANQJdHjzAQf7etsCHPJ6yZ5
zG1DQ2qmJXP9OgytlMAiTApfYCPS7visqoWxGpI9v7UHHj25glDsWtij13QLyJOrtQhfl1+PGwoc
0dgYFNul0wgR5/u6f57/s3z9qQEjx36KrE57fv3RqOqd90QMFZJBjiWOgFWZgsiHzjupImvl69/v
82FlRLN8eQ6IKsQASdJDI9TmHn8cO90Dmiu+zHani5FaMF+tIg6ZWOt4CgrkmruAyw4SJs1WBWu7
D2YWP+sMrW0g6QgMi3kLs3VR7y+DKQgqUmYjX/TP5Jm+ZuUrCu7Adad8v1Mqph2e8x3IZUlbs7oa
yzRBAHmJbeoS51tHEVFV1iMN5MIXX5bXnEjZ/Rq5ecLfFWvz9XHdH1fjp/cDWE8F9qJlCotmX9Rj
n1mmz35gUoxM4sBq5NlezdKaV1/v/ib9iaXU0NgBsb3DBHhCXyR9kW0uHNwAdvPN8wA3cS1ue/4U
z5oqsdG+3GRA1W720SbCEsHI80dfYvGrZirIE98SNHDOU7maRRXKDG4FVLcNc0BiNtewWhKtvlvb
F0dfbxVAsEHwGNSpItF2qlb43CqYS98Wze53nIwhzCRUGZfBf9zye1O5s1dUH3OYVcFvRJbKodjb
PkjmMLAL0EBm502iPUgLokdItaqo3baLRRQq7fAY23Tao8WOVevrEIlxEzffWyj0TnObohNIugz2
Pt7/gm6PoTZryqCK3juxM3x1Iifw087xUnC9eMMRpjqjqKXyiJeMN1NVronk1QiC1WrY+Q6Hja4S
+8h7EzZ1tFgdSl2zk0NyUuJYEV6Zx0CR4fCF/QlIIB5caCDwlKRF5XOWv8ocIe/OMhmatsUL10mx
WqhSyjAYaKW3iMOM+hPQQslzkKDRwHB+Jb3YWTZWcfQSnewMsKduND3IzxS7jrtRCCwz/O6lLqY8
SnafN7o+5o+XDBMQQ00GMw06Nrkq31p7yI5HyaUy/HKChHX5I1K3fg7mieR1OsIC4n5BtHtfkv+Q
L6ydNauEHwvWcX9moWW9/4PR91bmAUL/2ugtewPuTwOxwpOEh2LNlJkbvEeMxqBlMI1UNlqI1ImH
pwZKFMiRAxE8nqXzwl//jbkwdMRzOTHxPSxDNW5PMR2CF7TCP9UN0oO7yQVxDony1tm8VHkzHlfX
tYpIaAnUsv1D0/r8TVNwjh3PBcufX3RxkTUc3apbXZ1tagiGKdqOajlXkL3P0gK2yTIipyxu1ItI
rwYr3cFxE4QX0p93dW8bwUe3mAVzej7tIWFs2kC5Fe45NYj8As8CBExhjICZ/7B5fSpj8ZBQYXSf
bqeznE1smdRMVJx1cC1nq7A3CsTN2mHcMxABwNBkR/DztPwVis8ZVed2I9xX7aVREUuCFJNqDZIr
+oBSJKbd8dppkvJl2O/zLcGjQXz/at10PmXHA6cMOIlVAc4Ly8qmIv4Je2gvvNQObw5YHnC66MHk
2oMmLg6BXJk89GmcGlqdE48PiZ4IjKKkHTV3jb6P91Q2inT0dj6kkzTyI3tIxSBPJnr+Gen2attM
/hs/b4ixDDA/JbHiaRATPRhuIxwbiat7hqQC9alcLMaXd5jf4Tn160HAIBOHiGZAbU9Sa7F5Y3x1
sqZ3COWCsMnTX+oEsipfarx0ASt9a8PlLKDGBHf8zFBxSliKADVC/dR8vmVAqRf5yA70QI8vYBqJ
ZKa9MreyFowbVFvgONLWjlm25KEk1NGA7OQthkKAwln7X8ic2ot50G3J95cq3IBFaT2OvL1A/cqQ
xLbFwdp0NN+z4lF9vVs5exfJaeLoKEZBMh8oL2GMTIk/0Z7POwzKbso1ZfNFxmfG/5QAqWlqwesq
XgwArMNOWOodbZS6BN0gWL1DN4EhCQ01auViG7+MS8U9VcwhN1r57Zaua93eMfzHJpGgGAObCw4+
r6khSN7bb2aorZ5JsIOEeidZNmpk0hrWVo9cFxHY0umgOV4ref1ROjs5HEOGR7XtxhSqrrMuPTXO
ujFal7kUBNNMN7KdqFeqAHdfyZ8wMiAFCA93LyWxpEqNbbkPrydWkxkCSwvJ893P7DkMuY7+d4XD
NzVk4IRTyXU9ZBPmtaocMEvfDhx3LOEnTwbVLFCI5+602lN6K7VaPhNzM/MKFEvQjugKWPy9CMqA
PUgnH+PBy92M5kWvkWVasfi1TV2a8gBgbiSPFM52iAAaZHQ9xIRw/efnHAn+LddLKSgAvz1VOWA+
I9x3iw/5Yxio7bi8scAZPupQ0pNNsH84i4ECprctG3ShUVHysBuZOrKGRe3kVMA8o3L0R09DIYY7
nUcFfnN6D4fJhEEbSZR7OnbA60eKiXVIv64oyr64Eno6kwSPYFaXPpUhcY+Z780jvYnGvQKacHad
Cr7N+z7hGBp37TY0X2h0+MFxqt0gNkPRsIN+d69qlngQxBs3xJOCb+j9s3kJCrRzt9jxkj1TILww
qno8iet+pZibb62e/3EnNwahujK9SZc9yzhSiD1F2K9IdW+1FFNwalxqZgd9mGvUCTaoxYcaJ18w
0zJoMbNBrS7sYX/7hkzOO0ICEfNARZbr45byCBpyqueMLoD9y7yj9zhKMBs/R8H/WqzgRa9JoHEi
uNmnM/oF6/ztbjoZtAhvH8zijfm+/LFXf6kuVwqSdzZNx4x4NXimYqVPcvZohfBsBV0kGv/WoOG4
zM120vzGHPcpc1nWitkoGg+RnNaN2xpnfwdrfluEdD4DeLZ5Qngbs4JDjDQitaeV8Zd4mDEOE/Ef
HNe4E2rl14qqA+2mgaNNwKJTElyF6kPnOtCJ0m76I483z7LWhcID+vg26OC59Zje2QCHxtbAt4cs
WUySzhk/gYM/24e3irBvGzC5XdT/eH2oGyn/kiYJBCgb5/cl4JOBA13Ysydag5a8HkwCQ1OdX9P9
jVld1mNn79Xxqmdcb9rsn0L+Ksc91X//o9+HvdR5gDeIDCHp1K5/S83g/egvYjE/ShpgxNeKdZgN
skXOj7JjL5aEoNMa8Ey3trWDfTzoZtXT05ZBXlQB6wWUGct39TwHeE3aNrLmYcL2mSSwSqYMOG6x
7m6CveRG86Xl4AOnEnxPEB/1nIadVhsLZETO6WPPifvD6iVDoXSJRaCXk6VFXnsoKk+6ycRGOXZj
sRnwWIimHapRZRVnpYajuBH1p9BpvECLiv8h3rSvsQWbsfyUR+ynRz5KmJLa7AapwN051T/jNf7h
QqSZvMT1lJj/eOoL58gJdfuaSgWRa0cIqUNooqn2Wk4BSW2Lia6MEjTGJaVZGvzDpDzT0U5xhios
chLgExL8eTCqQiBGJ8kNNQauXhaKcga8FvmRnfjoQZvPTYnqq6X3RwGDvizCmuHVqOrLBuXUt7Un
Pv3oY0/+SYBk38J4K5Arytns+TWVq0/ky33mXY/2WIxit5+OISWv9jjgAh4gRGlYW95agyj8BvxI
l/Cf6TP/fw8buECw3tA9moJ/wxoF3THZwe5Pb+JHFLuzAvA+xhVLqoVXn9YQIWRcQJp17Jgnxebb
5pGJwBMNRbMmp6YbAp1dKRE3SUstzSLrnSvN2yHqUAhdDXsAS7GyscmyB73m5U5/DzCBhYvyEGhf
MNEuuKR2b4spS7XOIdEhRqIZqr1UVT54QVB3uBDSru2aWXweQkvOzytAr86KkBLdR0wNxuxR74qM
UyIEtJ7NFlcbRA3Bl9CtSOWRa6sPz/3Msw7MBEnpqrN7lMTrd36Jgsk0RZq11o1L/RIGLVSEpiD9
OgkBW9YdtqiqC06PNwnePdOxIZ655mDaC3AymmerXSDIfLKVj9odW446Wy2BshafNCWrkyKGEDVF
f8yK6xNx1mtOuMBC12SKH2Jd72PELp+7CNi+UVbryT7/iuF6CC5ciS9MXSv98HFjjZ7AKtmoKqOv
k33k0Me2+Dq7hm163QvGHTjSoDnidU4t5fCGhj5Jwf4AgYTr40+xfT/WkRL5EdL0C8PIDaM/tM/4
SQX6B0iPkaKYdZMRtmwSVEbmdZEpOTiqZ/GND2NOGRkIwVrCVbQ/5GTZEDAqpdrI+KZKNSBHQYVi
HgR1RRAeBvOKarPbR+xF3fFalHt+RSJuXNye5fWBYGkfxwvUoHzFMtxRifXJQF1T15gupj7TjH0t
NivGFLzr6ND2VC/jmR9BmnQTTejPcN7boo2to04yV9phnTQ58FKapHLWrUQOd51gcu2w0G+cLB/j
HBzi4zAcRzhIVlBubACyePQu4FchBmHC3IwSoqMGc2DPi+sCS+AbuZ6V80+JGXxaKjf/Pcg1UBwx
I0m4JWrbhSTuXeWbDs8RECNWohi5foRcpGxmyGOJ1iQUm6v0rUPO4Llrz479lD25q+NZRGcxYxFe
bGL46RYWqapyd2OcSY9YNd+R/zSpGxNLWhG/oz2ZtZcb/ll5KqLFeMLx1IYfCAz7ML7PmBeqqN0/
CbdzB07WFBRFzbDru2FFiKHa6zRS2F2wBME+3gjZKXxCwxcWqhtvTf2H/OhsRM1sFqjfzr5D4Ue4
kvZGaSFkwz95IcAwrF+HKcTJkbZObt6Rg1YVGVQ5yNRzgbuAGFB9PfJIehjC8WHrhm1R9P2k7OqF
sC6YvaUp0yLb7fyj3RNZ2WnneLSGyYcpfkF2dSukN5j47gOl3mpad1yLaWD9bhwjOjeM55Fsmvmc
8YgTjlKZrqNaHeVl0EjqvppQ4g2Lp42J6Hpl+Cdf5xTUkYAT/hw7SA4S/4zYJ8rjGpl/wd7Mnegz
I7/jMYVeD1mlUobm5VDkjNnIuGQv2RJFwGCXQ8BgwbLIvdTVN1+Ot22gV+pI4jvkcd/4lfIRe9Me
t1lPU/12HU7KJWvlvolbwaQDzumfmj7w/3zytMVCYAhQA0BaWQHIuZQ2I6gsbdQh/bXJIb5CYAWC
/1+WJmcycIIDrmKKuaBKO6XX2a4T84G16jG7O8LBFfaaQU4jbX+c5e+VNfX7rMKAh0Otd6szGadi
TJGSIEc1QnC9/oDbpopHGZcwPihdjecEb70eTDzhwc2RXCUPkuYzfs+zQz0Vmz35FoCBmw77DHv3
Og5OlLoriFysZ6AFJVtAFAnDJmrQB0voT7YeYKbzuxUjGqG7Hueyw5eqsI+cyUo3BkFtFuLi96Cp
hCIAWQFV7PIJMJId1j8WTAtcCL4AHQhjnW4Qx/2zvaT329EKo3r53ZCthLadcVxrcwQkehSSro1/
yWTZN3XF1LvMGXVDSwF5XHQosUltyuw/VsKGO87daSwGCLjf2PC7UZYG25C1DXVfn+xWLgfRNmof
PEG4h8B5Pku3DEY4OF7MObTVrF7keKGCmK0adUTfAYOQ+XAjKV/y1FE9fShoyEwAL2CXRxCEk8kL
3mfS5MvVwvGUItdoLGHcD2PDuws48C6aX1+2WtP4zBgp+zBaUaotlIiToOamZTOcH4w/5RUHUaCO
eGVnTvmZ6OyZa8O1EmrjsxrO01YkjIAMOZXki5zDZZf/N1uuGJkQIM29NW0V3QM5yUAzVj8IYAks
Ffq6/d9ZPTwePOvY9VBLXSk08/F2uYtBxHhd8FLMZVfebgAgxhqwa214iCA3j86ui6OoSwMFf9/Y
3ubwz5PMcAxJrHZx1ub73Is9UwoMIYlMNz3VcT3qfHcTlxuMth6I0Amr0zvu/iJCv7OLmxBo/ToF
InUp47C7MVU2K5DGKzDmtaJwa2OKkH4/KdfFlUHx6/5WS85ZgdRfCaurn51jjdHh7MfoozS+q2NC
PxFQy2NfifPjcfdogVqTg8CriOfeR6d27yI1GvMqwqLD7Hlir574Qhi/u4Hb5mjviIKQ6fwzPOiy
UzNTeJt/9kGHb042Q/LO3VtI1V/qHZah+IoXBBaGu+VPB88fLwN64XOQFcKTjNXKbL8ojbxjPbUQ
lw7ZYhe/akqM3062744yslbNOrdZRZDcCbJiHQSqWWXbcTJmgdJKmw8ewY2cUCZiE4UUcfTfDQgk
SMm2zkea/WsG4l4AmDKogCrTEOFSSXjyCNreziuvSAaBTnksY0eB5spJ5w0XRRFlKrKgQPPodfvU
fiqEYAZLrs+R12SzhofafW8FSzBa57AuzTk9jc44DoHJyz61Vja6KAWTGkhr2lOsy3UqcgGNpCif
NiVxGPw1SRe6iQf+7tQDL8jL/4MqXQTXtO7afoXCNcaAXOW1/RDnc5b30lftGudukdXImt93YoQj
o7DgEh8GT8jx6QOe2Y1myAvcRsxmO2jc2kgZxjG7wYzjwUoj8VhpBvqahOUg8uAmu9QhZjqgkJ3y
+cX3YLBxMi5cyk9/rMygPN5LO4VBAmWtWPQ3IhUJVQi6WxJC5DZHN64JX23GGElh0megYjMfVbqL
AHpd5kI0SRxDf+WfLu950WohnPZ5IHXVZpGEHoasacfPLcAcZ9fUYqGQ63Md6tfKKCmE/11COfy6
FO+5EcnRMyJrV+xabo94AZXKhfsuLliGqjcNdtPYLW4swwhJD186CyMbFEVcGFXdN5/UI6cEknzy
WCUG+C4NaAkX96VE2/JJ59/vICFACaAJW/K+sgBjsCxKg5xg+Dol1dA2hK0RsEwoV18e+z3Ynpgw
3804AsyyxBveZkEbmfqQx55V3abDrGGjS/6Cf9TdNnansBE1dWm0fDrLKd6Tev4H1nvi35WZYW0q
/dg/Sbm6jBC8iwuyCzsyJItRs/iL1BkUBa4B8dGIh5aN5HRPd6655MLXsXdncUtIMvujCj9uCZNv
khbBKmGRoB15vpB1pIfbB4EAtDaNIcriaPsoAQrsr8OZpxCUlSe3d8MImPMCQJTzC+WXxhp9Occh
N4xk6V9JhFXer4pumLDjH9o5+dD520pKhCzrEvTBsIOAFm5jatIS2Wr/67+wqdOpjmXrB1bFiEeb
GCicQ91c3YknR0WZkpAM+/rakOSJ92I1Mv/mlBKajJRybBc6oXfLMw6L3CfhGbSk/lf4znU9EMeh
0AeHmxp72JZxhJBP1fYJFF6Lt1zKI2hpKHA/VmUwzxWIalZ/Rc5u896NfwQKim3tjEJ7bogIVoYe
O4xExhjNvnUVj2Go92iLPaGqS1dpCp95wDrEMXVaLWlvv0/Fyn0sFyCHkDZMz2345Zdf5IsLjoP8
3dT5GyF8fCKg6cUSlBhqaidyHYVGoe8q0UhtaVSepdpiTFjUoye/MJ+fV/jHak9xaGFR4y2ZTT82
ZLKaRQ8bfmMbfxYbzKV8qbao+b6rccfWymARiLUCWN36u8fsWcN5J0nbndfrx9hI0axmijNed8bz
rGUB7A5DJQQNJlam0dlGhR1jMdW8gt3Dpsye3foB99VfnumTt/IQAYCOvARKr/yHqEeZJqOzm7DW
SM2ZPwbhZ5u/HChrLeDJzpmsoMbsRo3mjjJMYERlUBKKafsXafXmQOXK5tEzqAQR5HIzE0B663za
W4cWYVMJDNQfRfDF3aA4CaKg4WmFkger0TpoeJkD/ue7MXR8C8mGcZoDHZOwe0NQ/okhdvxV+vYN
GD11L7CB4X4HcMCA4DvZQBF4ScbfiWjTxM2OzfxgijqmwZDmXMpHB9UoUa4zyD4rdjXaJYgsM40j
yGkwosXERKVpoALriD+jHDgNy+CaGy4XlDPgblOEbu0m7WnqNMcrQpAypvD1bO+xrjajPXXcbFdr
LmevkxXl/ZLT+pbwPEQdKQEmlqEH+xnbXj8ralXvTvBD1GE3RkAFVU+K2q3oNO/2g5PcI0jZRxeY
ZUQFhYzZ8LXcT3TeBrvFvLwsnKZAHhbRZSXsTWSGj4tQeeMmDZu+Q2P5/A/VI5LhAF3/9qCwS4Xx
iB+yuqH1cVk9tfjsqkAfym5ZefD3h+9dGxCmuonok9uWIBHQ1KFjVhtMwBmgkda81lCInSmUe7sI
7wkepQR6sN+EumqWejUTzV/6OC/jTI9dQLZYVv8xHG27H0BlSs7S7n4MzQsRKGv1+Xfhwp3K0eCM
zh8NJYjmQvgboo/pPJsaukoYiXuzGhsaS6AiIve+733KoyBM9vsX6JLQSLBao2Vtzvmnk+exGwMd
RVpfLbLjYIKGwhc3IHbgo5Wnay80ESagMqgJE8VoXbVilbJuALH2u19QK+n2A02X9yJg0pEtg1Ay
ULj/9Jo9rTUAJX81Es1M/pfuZDAJnsenuh0SBwS8yPPKm4LKyBafY8FWfNxW73R2pGIg1wrQWxe1
OHbQErxD4YcoAI9FETEeE3WmsRInKIZVngJFSOwgMO8e2hc2IggsfcgVukG8Deegz0NXx9dngrXB
PoczP389Htw7ihTZa8Sf1IIBI1rWtr5SSlbDwJ5NS/TJji2KIWz0bTJQZqlCbubSMfDce0oSCFlU
YR0cpLs+V7DoTM6GapoNcAVyKE6xvKHzrOlD44OaD6E8+3ap8aO2LUYeSHCdddv15tPRhgUxaTnU
P3aphqRbiqoaQsMbNwlYGoFWzz3DTGRri2zw2lyoaAbjstjaiZCls/mYhfUlFNVH55vzkgDpcM0g
NoObydqcyF7firhPEL+kkb4a3wbULIxeDtohGvpZmLg2nJ6DrwqmaEgzgiRNzd25srB9koMwXcGV
ftoOk5hsoqBtioSIKRrXDs9NkQdgNBzFv11DbQHKBHGqWSIXznmhMlRUDdNUTcgxedAncSXHgZGl
QtJhSpESVCixf60+rXVISuZS7xoUBIsIes9uxTsVJeE7/RpX5ovVLqyNW2I13HzBqjz5xCWqPx1p
r8GBe3B+W1gWi6NloNy3a1HxWRDsnhEfNTySoLBaLYPYcbIy9G/uj8bwP49jzeBgW/5NL8rgUq5B
l9Pk0CCbNTjyTsCuUwfj3/UP8CEL4J8VhioQrw+Fu5VA6jUaN144wa0l7paqXDbdidX+CY8toRKi
VmbWGNPGv5zjcawmXzYtNW+BxnFz6pIdP5vBcte8k0B1Lvz6yDXZ315ok7gcfSwjTkrDaNiFVFFB
ygnS9OJ1EawG4mzbIdxV2feObVbv30rASkapYg5JvAJLThxVghgRdv3mlowvGa2F7UVD81ZtTYNh
8D2JuluYbMMH6CmEDGgFf/b63vg8sZ1TMEdzOGYj51UMyAo2NUndh8tWzUWekPBc6qtLnacmfmpw
pG38a09GzcjtracaqMHKpx3N4Y+AUafgYDTpSzFC8SCyweTw4sqdnBC9JECkRx2SeDk4z00C1i/A
PmDOZ7w5qRMhjmyFEDnI0PjdwIulxw2VXe6VDJEhhaiB+YriwPtC99jFi0aZdE0d8XDF0yOmfMEl
vMxuegaX0AkndLmerNNA8Lrvkl8A8FWfdp+hY6yG8tHgrkPcP5bP1xYLu2Ks8TNAk62xKuEN8E4U
lTKrlRoC/5M0y37cM0vfRrGrEJM6e7bYpqR+vj7qIzVXSGC2+8xDV5Tqmt6NhZtnRCf+QJ1RVVst
kxcpWWIiNFVjA0/Qzt93cbzrKEJ8lXhcrMrTHPA9qU2+ueNr8Y0yEdoKQVcGVKWPnfnYiVhLkwko
C8DAinZoy0aSo86bULbY4pxcRYFYZpLCE7lUSjvSeO446hTX/X345m8+jFscw7RtFYNUHh13xn0F
40vyNG4b2bxZUjlrC6AG5lOI/LPfb3nCxMcA1v+3cWpXhZ8eqsOEc07b650myU6qBoqABOFiCZNw
3BmorM9nw04GbdRrPdgwGd+saUQ52XAxQyRnIqkRR6qoZs8DpJzYpPEmAaEdRLgWQfFEVR/EiWcX
Lw2nnFoms+iIio+hE311M4vYfVk/2xOfjwe9BIJZHGSKNkqrK8G760qdP4SYLbStO869NpVV1OOf
XVDAzDgouIlWUqmaoG3f0NdIzci6C/xFl7ylFCli9iPCJn1oeoIzYzRrcJGyU9HDvlub7HPP7YS9
h54txhSplgWW7BGCi2oAKAu4PqQnC2UT44tC2NwK/U8J813FRTIpa+WImAyyvO3HJsRO8kPz1O4P
jQ0xWhXC918TH1YouQ/xmAomYHAMSMLMff1mOmfDfvAHPgVJSzTjg+vpAcxz5GkuLUOZ7JMueSc8
CyT6H2sW/J3wYDS2UxdTX+gzTK8w1UyFYW2zGGpr4f2ERjBm+WYJc01UopKst24giHVJAOUwfgnK
oqdXdVIpRS1qnmO/rQfR8Og+94XOuhGgFHgQjGFwyPSUC/D6J5cAgPSo5m7/uHz8AeUhWyuWChFr
8oYFi7OePq+SVvVAcygtUOl7yoOBum4Np3EOr3Ss3CyCDQwQ+nO2xcbc0Pt9w8yuMOxEE4t73ypF
dQAkra3ccgOMkrYOF6JAC31rQv2nTT5Jr9qqzm8sVOe3ivPb108crtdIkWv29beGQjiI+HyNM0ee
+Ni3KA+0eGUYHY+XRTrsxUO347kga+tERfd07CNcgjquVuL4wFZGQ9sploVe7dZ3YiMlaCe+ANOG
36aFy3M4iKH93H9kPlnRhujJgbYyH9Nb30Dsw03WeZZEe5iReuQYDOW0gOw5SnFSOwapGmAMZQsn
EWdGq84z++127JigoXiUZl4RXqWfMRTVPLQVyeRbmL6QXDtXPN4pY7MSM0kh2s7NWfRIz7WnMIzD
QfQKpvI2U15InKa0tMgwhV8m5opZWwQw8KrtDjpzlkE9SCK/AGy1OoCaL5Pbp/bpDr1Up913QQrL
wO8SWwve3DkH2cg2HQqjJ1V62MUBVftQfCUlldmhGI0gyzzlgieNuP1rB/BcDa1T696aGiNwGVA6
HNxFwy2OS1ZdtZSIBfGoKMcffaVqTxU7qDLm7OrL0eYQI1bZvzJfaiqjcnzLqZ4U1xQqe+VO8k3O
WWKUAPqexHVRG+85Tl4kR5AVusOB/5RrjnjpVBLARDrXBLi3NU84XAVLeSAmiBrXLigbm5jVUFJW
uu0jQjE+KLjCrsiG3Ya8m/I/P0+YyLAqBpNgBD62OMF6tzKHyhmHlcf2O6plxdijAN+5mVTx6hrm
I8hH2yyDfswg+6FULTlb2yVyFJuXeaxSR8L5lXYyq3KLnzdyc1b7iMLLeZPClxcYBXu00EW7Th2T
iUUMzvx+OM9OmxpecMK4Hlbg8IIt8ZTQnJswGsr7FNOJTP9x5ql6lG73MGwChQbGIRqUaZn2rwcj
8+EYBgr8ccvkH65ODuVoFCJRPEIpCgy+9lQv6ExCArnlnD0ZaNxnvvi8F0xN+5VM32J0CNYoilzT
oXbhhnlV1aynU5geglsxxRuThqTYVqFUCHFiKs307DBGhq8/623B2IpuUUkL6kUFJd1n8/VJc09T
0i0wCLfE/JV5BK7E11r3d+RF0C1Eg3O/3zldr7rpMy1J7njRFyoIDRdmp1YjvZaDaINXLeYpBKUG
6uwORXLVOdQ9PN1WAT1xy4LgwI6rOiZK+R04S2VVeUw8CZNp9O6SNE8Dm73gr6EeQqxI2OsNKEd6
Jv2xBW5WMl/G2vyFezWKJvu+Zu34VzsuiPRLM2azo4E1bZavOP8M/L6sZylDDDhRzOxiD55B1ep5
mhRMhAJauZullg1Wrj4jPukyitilnU4HkFElTViBbu1kEveE0saKeD0efV62xHBba5zOjJzNqYfQ
EZV2Witc/Fy8B05AikaF22ReUD+/16ojjIp8LAkj1kvyoumCAIz0teq05IiBHEexQmoSlPuQOl/Q
UXjLzoPZL+VAx0nfb64e3DgmBwSfbv+Bh4JlV7X6bFw7oPmIPsTqRwamAY++/BZyVJVtRLxhh8np
oUKVgqUwUtws9RiqNzZ25CTuP5c4/QIk3gpAZWITyu1avbZF2Dw4i8kxOx1LEBvGF1WpYiNoKxrE
EUk491JLLL8zv5M5nXz8CBTZIsPfDq0rKOs22diPt+MtC6zgNx4hIwh4hKQxtC9Wxo0exevD2zcA
p0exgqvQ372lYKUqH+q/i4PNl0dnanqtzvcKoIpywOyINPwTVt6j31eRYb3dMGtemgaT8KveGvYM
sBh9iRLc5zRdHPWlEnG13Z6rgXkbSS4iP0sOduAoMwzo+vjiJDVyrRcaM5jSYgRnqkdPy+PL03Ao
qwSRyP3VKw2vMmGBFhbKZwMcfqWXiVO+z9Hj8bsR7c/FdjrTiDSMiGVq4EJIR+lJUvcqwILqwgNe
s/9CQzJwAwb7QjcDIPzmOJ09Ac0OwgrRq8bfD15bToeJZ9yN6F+i64QREn/AW0vWorRce2zUmrBt
oe+H5uaAfxq5e0u0l7PBW/FeeP8cUohflZi9jvZBe0KIm4zOSZOQk7j2cR/8B2oUUuhxM6zXkBBd
tpMeScEQG/pES883T3LYV9l9aATWAOjL4PboeTDxBqktL+qc4kIshFAOENLzLkp7gc7TE6d5xkjV
hSdEU4VWZG4qHslaO2Z3RkuUXUHVSGak0ZM0fI50Ju94i9qqs+BmiojuuWeeKcxz1hjAsQh4lpaR
vreTe4vWHkpZPn7hj9Z6UtC3wmSaS2cKIqhYIIS8OZ7ztqohX0ZQsgXcHw4k1ghFVCd+GL8SJcyE
jMHwFXLxZSR7b9svP/mmzTXHvR2iy6q/PyyGvFftDDROMDQSxY5a18uW/qAR+MheQ2gFzojlxXND
e9hnAVhNfrrytqX8MC3/h28d235ntm9JLmti65MqemmEPcoFcOLDx5RzHUJB2ii2mpurOhVWVN/B
kufUbdz0MCIFY/jxHFjVzfi62sdx1aAlB7390Uon+Ow0AlrtI4RhbdybAAMtqW89z5VaHun90Doj
+2tFR+z4eRwqyWJu+tSxvU+BvTQvm3RfUhlLfcVRZ1WUHn8VnO8cwNOGy/aVyMAeasasWsigDmXa
Y0E7mAmsJVIK5upQE5WemBEHkMvovo9M5+oiMeKYjmJmQ/XeEZ1ZwDcETkkPMWlZ+5lhy1RQUSCB
nQ2VQsE37DbjxY5yVxuGnctwYuj8YY32GjOD8WfsNjtB1Mq6zAJZtNbS7D/n5C7+/ssOdcyiZ+m8
mznoSxM13RAG/1alOLsrK/UVZ6XzZrqFTqx4jZOWxnwpUgZxh+G8fUEHgZ2cQTg4549b4TbNqpk7
i4haKG9Zx/tqkiYa0Pto9r+ZLNnE+K4gOszFubg4LbF9Q4Y/GmUF0crspoFC3bwtSBE4JRywc+/p
ENIzI3JnPmjvLdd1dO9AUGTciwtczx9XSTrL+P6sKZVzfE2jT+NyQRQbrCRzcaWXRV+w6n5+zghf
qhGV5r8lVRlaRrpH+RPENSL0k5YSOUJ5N8PNr6MbEBtyebUSXQgWlDBOvgI0tBbAGWpKpVbvKJAO
PHx08X0PPJlVQlkMMDi9jgpNmOjADKoxi835p2VnIp+EvfctQB7Xw9OC8QQiTfdAM5PeSRsbL7lO
NUvVqlsYHudk5MLoDVZted17XBuU8gIkoGCdlUasgTwFbQ73LASC/CDgv+hFtuYWJbllXYQPM5sM
zgYLAjmHTvuwupdSzmQQiOL8z9NYG8l7mcjnyrYtVaMPtHbx4bNN4yRJ8yz3GFQNm8XK0oN4lz/1
Jf0lvXhB4nGAKNwkY/sJocupxIpOeyOl2KlB0/U16ttBkAWKYqDqEvndR+khO1qoMUji2LdgZAlN
p3SD7TttBkXFZLn+f+gnMVCopOTglHb2toM1LSAe7p8mRx1xQkJ3wAQCXXlE5hI5SKM1GcnK9e2b
1BOVmAB/uEAkt2RYYYszsX9hmX3Ibnw5Gc8FS8j8sIMBsZOU3bGQb2y9tyGFsXU6SuK+Zacq0CMi
CrO8KLW0QzNoUumKF7+7+5ASE+B46x96NLMBcYmf6auBgHmOYE5Hof/VQjTspRGLttwbRbrXgcIr
KVvhk/qsAVZacJbHf/KtqiR/CzPaIy5RmCjno/1C50//HAdlKyHC6OdK2F9SL9Cycsk9gkq2H2SQ
IWvSRYIAxNT/TY++zGlpwwKOAuSboZQylfMVtHnIGx2OYHHWam+Xx7TI7mwVqCf7sxr+f3eAY8h/
3A+2Ttile9XQiy4AqOCa7UrLaXRG/YKV+CvaKfUeNiHA60wFxPQC26drdUcdhEmSu/5CPcpI6wHl
yke2SrP9hoHx/YAWJ8lVZM3UCqT/8I9FODANoufGNJjKvjgOGYXnOanQq61jh9APheUqJIyuki6l
yerf/kiLIBMksgVMH/WYROfS5n1fPVDJwCM1SGXGPXEhL8Q4IjA4NFCShNcMOUPcQFzacVUF3GtL
5wR2gymnKxozG1Md6/OO7foyHX+tIQJdQR6YXnLGSEP2vD12EMCDGaHjkP1hc5+VT6Kysv1dyZgX
pBaOjsAqjjk7Upp+HAf0KU1b0S54lcjA17udGuyNheTQU2B0VlFu8h0B+v/oDdD0hxZXHmOyKrm/
CpCueQEkEapD0J8AD07LQwUYidRrz5rQ8kOxU/Fc38qFt1Y9BEefyyPhRJhzClVEbyYhA55OWrFF
ZAeMDLznwLYvOhK/uHuxBfuLcKBWueKTsaHwWUPquj2RmGTB8nO1jaCFf2D0P5gmdBzQ90TK9wAm
vNRpFL38iEPIwAhtNXZMndBfICQp21BGVBcTbreAPtHAR5Qux4MYDn49xaFuxrv44cMOG5FLKaM0
1F7yvtwf1dPISBmOxTsFETxwFxDrNbI0qZAqIGKYHzUWRmDKft1V85fH9fblDuAhgpsIoz0r4V/R
Qx504Vk994kW7ll+azJTSBsEjtiszNvSBKJC4IHg1FidXSYzgfX6L3OjydDauNdYNGv7ntJ1TpvA
Ei/NdqO68HcpfpfF/SsZjDJNaLs70cm/0TaJG+v5Boau3Ff7VwyxkcW+tLte+AShvA/xSxlSWm9r
wgrOWtSPxozJtN2543tmVV/IaD869QmzJrFjme5wQKPUT2LksHMJa/bStNyLukanSwmYx1zn1OYk
tkO1sbPxPl4bIjkDJ72yVsWVcY8lNhIyGB2TqxgiMik7WGQgLb4vbyGOH7oFS+y2CL9b7xvOJhkt
Tq3KDOjNJU4ajCHfoKRu4OGjiS2pksck6xs9ur4Ig4KLK5MpzrJIYqtgrR4EcvZTDGvX2p4chYo9
P69FfIyz5reXn1vWzBwrVC7bsbNoph519DcRUmJi8rcFmaUuj/lATJ3BRNnAHpch92aEycs5ljHv
/my+AsTPwJebhzrQUxA2gRQaRTu2iRfHPTpg/xnqyBkxg22tQoV5Xttd7aMcsfd3LnUXyM/lB3dl
mMym1sQG5SbGisMvjmGanqSi1hXEwzeWiTB5pSAu7R2gKhIb+kbFVFaxi63S5PeUQVH8gudNkp5v
tSPtuYlY44n1nEjnjdpnYmnjlbg2ZUUlYjHcbURQl+Ov70P/wxpkbdlxsw2ddbk91lmCJQaR5zks
4zRFttJSW+p1k9NgdZQIt3GZSrbc8beBKZt6opjJyyL7OgxmdvZmUY2tYR6v9w5CvAEnktTY2vC8
a2uFkZxCq0Jk/yFwSkn92gA0B5YWsDe116K46gWdy/pu/LaARRa/BXLHKdeP+Gsm3xBmg2bNcR50
BAaLLkIUpTT+EgDVVtiAt73mP3menPRJnWbOFid0Vg5JzeQtqxpYtWH0KSqFhMYdh8ffGXJShKz4
fDjENErvE7oPeM5dZbBw8wmZ7v3dKse9irg1P6bYpQau854etIT5/5dY+L+LHRw7C0q2nQEw2BQX
z8TFp6oD1WGFhwxnlPDYVhEu8iAvG7rsxbmFAmhNY/8S0KCXr2Ethn7Rbcw8sEMT76bZYOwg41CE
o0Gmm/5B+fuTRWqDR/XfgOx8OSLnfXnY+S8YR4cl8gbODi2uQU61Zkv9s34GbXVcPehGUEc5WD59
Aa7Jrs23IWOP4jx092HU+t29JVEurMuf4/wp8zrEMN75/dscWCpbJy+gWOR9OuSSZKBUtZSSUHjr
Bhe9FHPPCdi0EHIylJw7jzqkTI8nM6eqWx4h6WmUZ5v1kgEhlNyQGCEDBPWOI0BkfuBhAjwX1TyN
dWFQK7iOhAdWKqbi45/p8sZ+DWuuCvWOpHOZH/fDEaqSnM+/xfxQI98DEcvhqdhpK89lndTUbcb5
wswqpreJDdClcCyZnvUFDegNFqJ9Ge6hJJNa3L+bF6ePBcrYJUse6UbexmIEO4G3ILDNDJpVcTC+
NFNStvpDo5qI9ggPrCmEiVcrplz+SMBQbFJvP1Xfl9GzPVCCaeNdeTcqA0LryG+HexFOx5Ux19LJ
VveV3lxqkkt4QHkp4cBgL70/h0NdcwgMBVbfbbA3/WTiip5Dt02XJtdCjsaMuXcxbVkFbXPwehuB
zqwUgXZ+LersFXNLI2ybLK4/OqgXdT4Lnh6eJVsY9RYVdftPGY//+Bcwa4ALd/BbKu53t8ybtij7
IGRBfwTao/mtnoVONwcj2q/ZYI/53Sfl1mYUNsrmJr1y9UQ7thF9+ffnmCla0sPNUky14IaiAyF0
jgpXTuj6NQ3lOAzRAp9fqIMoKL6N76GCMgVDG9mrOUXI3eYOHFkr8sqNAcfD6GVdWngq/M7u+NUk
QtSWK55p3j7d/FH8rJKo0kx+XmCDZ3vLVXmOou/4fZ5Z800vzDp1oQhnmVmNx9ziBfRSpRe+gCVm
FqlHmz5cleugIeqrfENkdMKOUKpLyIXgB7DI1AI9ZlkxRt3mWWNq3n9JKvHkcWcdkCkVnUmJyS8m
bg7yktX9iDI08QmhivBZZCIJbocDA2FjXa0b/ddeM5tq/NW0SmxewHvO2NjIk7v5PvVBXen9n0Hf
b/Y7R6PuAbEFrr5aE6uqpuV9M0q9iTXrG5v66CVcr++ucoGqBzMXUOvIdVylSTFbeSzZuzm4wLMI
oOMkzNJJ+MSQHJfWwZ5kv0lZmJSxPxBPrVNB/NCqI0z1aUaR7ZzgqGCscrWaAA+WidXPxAEkM4E7
tAZzbt6Cy9CTeZGMcSkHSXaQcRnT9wRe+JEyGy9yU4Nq9yQGCy+X9VyKap/E45WZeQ4Kwj9OqXiZ
+qmjDjjKZIu+Iu1roIQUXF3v0FFv9WjmlgkSoBz8aaizs6TVw9wPiH/zYJl0oUOXbPiaEHiMpP7Y
x4trW+CUk/q84x9P+uXH35pX+GgAfrIjGW5iHbY3oat4YPltSOSQQ7v7nQWnWCo/CbH8SbV6e5XE
1B2n0bbpGpoH47F6nZ8NdZ7ARGE8hWqp8ArfzMLF6ytyh1KM0sEOcvkhAgHQGa1bfFfp9aFHR5H/
AypfDFXpp33IVgYD/Fh9Ysl9ozQ/NEt8el1YP1jtKgEPcCgMwVqPeO0z1/ooLDb0OWyHN2JhzmeO
4kJs/RlY17y72XUgJ5Q+PN97fY6NShkm1WAMlT3f8KHSf8cYxL2KZyS+d7Uk9tx0/H1O77teXEje
suZ6JtkzUk5zTLVUqHcLg0jGdnVw1lynK0GBstBvRz0B+LCnHxRkrKT+40o9ee5M2Tk+cvWaFDS4
tVN3ts2PrT4R+sL3BKAdLcV/eVzeVMHjWX6DZOCuiczIvsCxOr5Svr6Bw4B7BgM03UciJwqne7bb
7Mx48RnO7/xa7BuREA3nl77DNe2RkTYqzO9+uZU/JY98PM/Ee1qsS4ginRoHfuddVmklzP/ROS0n
8XYQ/EE/u8F9xsO3vt5J0qzuHrpKeQ8EA2UUSCwt2tJpcR52AwqIT6tztQnBCTMLEcTX2M/i13hX
H88HJF3XSJxFV+ttSf9FlY7XaU33C9+2MXItlKYgTKQO0idoiSvHV3Gr52cMcMeqTXc5yiqjlwUc
/qgI1zJyeDx0sv64209wDRuN0m+nB0CvhkQep8s1pRqcrQ1keYUqMvdshmZ+CuXhD7QziefLCx75
usSQ8EunIsl/YNxfXQboAVgZmqS6OhykSAmR+Wnj7Cu+2iwSxNvV+aq/+NSpMMDQ07hABF8w10Hr
UOz4NskWMwxgzHEBY7MIiV1OZJViCOGaytmyUgWbTcXxmsip9evqjYfbpPW+F01WxGorclL3OcMp
HhklWLe7Pu1JG2kCuA6+5/QIzuk3xGN5wo78eEftdOYLugcmOyVvRtpnTVOEqjZZaoAhETowvt+i
r5uuUjvDNvt1mbWjQdpEnvRaBzw5dNoU4inwmF3/rxq8xHq0mR/UGRKtuWZyK3rVM7Ed4c+tjkmt
gzJpssL+kIwAU668Q5gr0yFEKDRktEUGhAdmhVN/E9efJTJHkQPV6HFHtuqUn0R+7uXS+Y8/JsYM
+aHh7BvV0Vm4LXj9WVF8yme3dXrnpB3+6yC1IJPxepOIhFteBsKBKOPbxVISdpELFeBDcHZ5yJ6c
VNSQcM5WSSF+ttlLajkcpP3CLOEc686XB96nq6LUlRi73wI+aDhmxE1NcvmJOLuVMQm9KbEBkr+2
Eix1rqwoOWX3FTX0WfYTPCx/is78iliGioKJ4U+hNG/XOhHWLPPBGdXL3hNTwHYJ+By5MUEll++H
IIMUYmDZCQexf7o7qwEeCEkMgQLB2eIldp5AjeORW2aCoHYgo4VEVDW248VolPm+L+WKqs2/wmZw
+dfgqRUayOPfdHHP173ewVEztGrikarOe1Kg6hEEbyWFLoZIt5lWc4e5tyQGptmuCh+py7d2JPH8
cJVb2G2u5LSLVzXXvqdjNwtz86avtRQ7MdenO5zL802pZKE15Gso43PjzzTQSdPvJuzh8HOqsI2Y
yT1VlCIbAIKwn2OIvbrefVY1vcgseugggOHHVAcWwhnL0V6HZGPnVvTpviAJvzRgc4HLXT+aX92O
/r5402KqyhPmh1HbQMWQL4uULlrM5SN5g2X5mZL773/I3Ld3Z2NG5bvx0fLEP1NFcun01oPS3pqT
xmHegvX0raSfYBKjUdLWkLMN5Ts+CiV58YG1jNFrirDSdRq92FHdDx8aQZKfQhGtzGg/jb2EQoHh
V7poASs5/3DB2cDnjr1YEfD8k81noNbbB6HtZO/qWZpumbepwk6XYGJG1YA8HX6QKPqrJHm8kurx
V8Pxe+m/LeZ4FHG5MoTEIlOKs1wdlh7rQ7WGHAn2csEYfRkUyir/v/SMxdpiw9Fr8psIjtJmmJeD
vKe2XZYl6ZBgVh53Z+tmXuqtg4s4iOxNTNdE+IfKc1HkWPwPgQJNikYHXfPOP737PinUxu99o/Xc
ZhtJz/OsNntGSRygsGvV5BCTVpZHIqynhr3aqMrBqVDNUgzkZ923CXI7CPuUBPBTUll1dqs9Irfd
BvtQwzI87xn6Ys1oMZL6sW1+7/qmG6kFHwDORZO6kopVZM57SYAD9x0DEvwJcYCQFBy/Y85N/5OP
EZREZSYdxmAmftcqblVh1QwDxg5tQIJ5QZR8tpWvfcGhw+GAgKbCBOoluVn1ckcgSSNEnjOcQDgZ
AlWUh/augAt2gv7CkOU+4F88H33kHdeeCF3FmrJ44pvKCqqQUoYj9dFArHh/1iISsOQghCeuBjxG
1mV/LGutl0bA7jrHAzlDIrFqQkfIO5WutkOvG4R16ZruqBDRfyNOQrMINdCwcQObmbZUbOkjE08F
GDY88uK/xHp6IktZmx4uLhNHyjbbf31h9pC4YwZwKg8dW3spZkKwrCnV6IsRa/Y9Esf8fFzu5HL6
+VcSatbu7MBJIOBKIReGGW4Hr9ziAeK8nclduJp0R2emJ5Q6z8tEWyEzkvOPO8s4SgYvXlm3hvi3
h3Gyscjfc9wG/QHhklGY69OvsT49TYRkYHMh1aAAkKzOCzvdZFzeghMeoqclrnr2fXFTHvBmcDGD
VvUgCw5rNWOnfB6uHX5bamncsfdz+lFFVnv82fwmMxP7FsO6G1rhBansxOY3qoD+xb9QSSW2wo8b
o+fS5Dy7xUJ8vYPKUJYy1l7HH7agtmlsgHE0gmnxWdVIl2ExJ3ygN+ydF/5ICuBCQ2KJGHKDaiAL
/3y5E497Xw2HsPZgCc/Aj91mkWusZLgidrv8AnrIoW/Q5pFRu5bYuH3MS/WlMI6EwDAvvQVcsM/A
XlHXjgoqgiZDd24VSFH/T481/dYOPutooQap/dEoEfS+jdNA+eS4WH4+KlUAcvr5vbNnOSJZLR0w
TrOnpJ71Qp4SQHV4sd+p+SKEMhpldcS1tw9b9bSLHpQ2H6gq2P0h0xInOLxLtjDwH3CTQVUK3SXJ
4klQDartzUMCZ8NQJ1OsMv3ty5AAgHxKgdvf+D4CF76dPch3aX0pwoNz/oTEwIFX76rhR6tVbS7G
hj/CojMEkoPjlTI9agXVX6UpJYSpFbd1VFfQPnstJvzfxCwXKuQthdATkaMXvctA8pZ+0FuiCg1+
aihaKyel7j1CY1gKAtGLMVBtLxbSYPMBW27QMebb7KA/TTJFs8LM0Xf3GAfXUccWQdbpFzTs+PuF
AM3yHcVCRz4BGitNjW22KybXQ/xFWDItbnsIAn0CIZERhQQSPleQD5zJuLPPbAK3jBHm6J61IK4d
hv97GLWlE3ph8KKhJ6Krfy73cccxa8YiF1aEkx8aiNLiGarQK3aGaX73dcIqM6oPO3Foq9fkYoAJ
tm+rjKRqyPiS1TWHEchiwBCZ7kA68QR+N4vSNsaWux1+59PzQt46ggUe8Wz5JMFrg7wf72vF5ckL
0WvGthAI+S+RHgsAemiUQhcMpDQCP9gKnl+IV3duTgKkEsUdrGvlJO41H0SGDKv1LJ9GBA0SB2AT
EmjV3HAif+GLmKk39ojXjNx2UhGod1tcmkqacR2ECKm0ILSazLHa0ZJW/NbP3eZUcKy0rmlQs6iR
+hOfIFi3W83lFiciL5aE2Vg7nsU+jj2B2r52vtqYBHdVDlfOyfk2vwIdXy47FNVp07B9yUOfmr80
In6fumhuht3UTIanY/7Ml1Qpt1uCOBxz81mbznGyqOgpQg+RkZQ6gZh07LOhnfF5IrbxRaFaBhti
5m3J7K4M+SAiN0hoqk3cgaOnqAvMT6Fz5iRl46zUB1Ez5saYEFuHX/yGbcso35jWYncwzH49ZdNN
txmHfQNYPUk6VgAZHDjs2TaTG4VuqbGbBupzw54U1CYco1PKmEbiJZ4tmUyc5Bbu/WOfnDuFfqmH
6qFuURXQmkKrExhJWY2bjy7iXjHzZ51sKzECOLZNAhAXd/q3f1xPifS7dDqBNJmmxdhs5lSvjeeo
IfOppsXKA+twnFfvHPx14usk+ZSchxhlGauNTqR73BgbqIg7dElsgJvbdZVY2gSFsRR8eoXnAfUT
Nlu/EstjHJFkTZ5Iz8juotbWTF4sw0ixMOY4tTWDTjEd6B4puuEqtXXeQAV5ztF7y+mGGX7Roqjl
2WbCTekHgtkBeaBptHv6sus/8tGvnH2CcUmtWdVnwyAQzGkmWI5H67tM6hpKLSL9v641Mrz7JZM4
1Td7FF9VQBiw+/cazEXgPRRdwp7QH9zzyt5lvvW8KFX1UjAFXZm1lWJSGpKBT7HWAjrZgAwKYBR9
iWOTse3LNqSDndi/gL8o0BGhRn8za85xP1JlZhsoO0bAp+UwLddG7iH9aQAKhPAX/qLQtHsdf98U
CtlCz4rLqO8etULzxPM9rjlB8UIh+4SriRT3y/GbJMIjt0k4iQUNoQyb3t5Aq3Kx/rBa9BuScExm
iriYqCPUBzDkEQHrCsqN+GAYM726BCCbPHKN5+YYS7wDjiNkbv7wK8fqt9CIA3TQMv0mcShyjC+T
+5tuVvcLgC5GTKw/q9XYdicGc9Q+yCBWgk8UeQFsv0PM0pnxI0wXBb1DqMwCZIR/5jjwHZJaOS8L
ESlrIORMOJWPSoX3LNNe5lSzzX5fg/QcN147vYoc64OtGdfx/sxZ3MFE3V9G+pb2I0eMvC4N/jSA
PS2/fkLHjJ2eXZAGKdRnmpAO1oqm2ltmyOjQkudZj2je2WyZ2i473aO9wJ84ah43SEwe3ABO8l+Q
fgEzE031VDGn7hT2fj1kSbBXHrfQkInPCWBDgxtcNrvn35qNklRlmFuW5WgpN5PpH1mkL3bHj4S9
4+1fEbFHMyxpnPflFHy4L2m+AV81uARoCUkckoGdtirkwfrNr4PKoWTFa7GKdOfcoZsNsrkOdHNN
aopSCB/qm21CYNKsAfPZRTwd9DqHAz/0qEL2KSZ9Yw3hw7irWNbzB4j78i1BGQbrCi7LIF7QBuq1
UjURruOOixaFouLhwchtcRhv2yM8eWBJU0X8MFW12pk8InoB7IEXBbRfgFylD8uTwBEioyuFjeC4
a0TqQhXOAganErRy42Pnbxo8UMux97Negm08bqrkpUECvalnUIZzYm2Qnnpv2CSFAZLCTUOGKemt
xj86GNLbK4xabCHtKfDr3HSkDe7HGMmV9EOjGVidZVY+ERJ4ffrKn4sUbWgIhCsiIoQJVylpszDm
dVKeNDsFW8oU6Zx0xiIQcShVDaT8qnx6OFSkQc/SHDReMtjZyCfMtZbCVN0fRkg7ZsL0H9MbW09l
PDWmoZi32XwzVpW6eevjcta23JAKLkZpyN4iA4WD5mc+s6SS+2qIAW4fp8EIWeDVWZ6pL2paEjQa
E5n4ALC2S9tCsQb2NYfFeBAe4eprKiL7rLub5UG7Qbf+Aqd2XSXdRncKZnBlG7N6K6/PFkkBKBl9
UYmxeK2vu5RCN3IW+95EEXWjQxPGQPOsdj8M6RIdhV1y0IC7Y21YyTYBklf0d1N7des6tLcVIlv5
ANyJip2BanESCxIyHotGxu5jV7UtXp2XZsbKonU4SmSASHk7KHP1wCe5VTQ8OhNuKmJtF7t0ftow
/cnz6EYXnIvbwXUtC9t3k8NB/bGOo0wy2K/MSipP3kRujJhpZFGjfrsWQqlRx/R4EUje68NHdJ34
fSumhk9b+JFm0NC2IUgAzh1Nt4F3MhGK0fYIcj3mZuqj42Ck28r72peimq3/GU96xxzOk3SS6RrE
phwkFZkmqU2bFu2dUft0mdycuM0+WcX3IEwFQFygSnJY/vCbNB38NbYl0w6pXh60wNPM20n8eK1X
5Ig0yvR3UhpME2Cx5jJp7ITkkxkwuF8P4fCuaMBEnBEnao8FG0hlYRSH+6IQLiG3trJTZzZzhLHl
qQw4OMID+ld+44n/FkU3ghsMvLlAcmhlF01b4q444U9rfl+XchXn1Ksue6y4zOoi+OBI/Rk3q/vU
NkYRhQMrp5xw3UdvXZLqvi4dK2+5qUXO5bvCUNqzlhqQ7bsj/w8rlJTnGkoGmuCG6JgvhM9hReuY
NBGI/ubSdFdp3NXyiNEyqGYadVVuVgMsiHWABgNVrKL2IL3I3CGdPla6eJym68MS8Mrehg5UlDHS
N8Z+5J/HXVkzAGGFrQUYpgsrPtqCm3uwGEkVOr5DeF5kdbye0CR5kJzhmfnj4RKeHHGLA3RNGEcL
xJ2qBiNh9sMqNyvw4iCjf7GRannK3+vAQKe21lk6sE3cQiQAz7o6YtpEJ0qF6Cab+IpKlfQOhfJg
2NkjgsGHDADE/nrDFunxpjkWC9xQpB2IB5S0JrHghDiOuoHVyIb8nVhxD6oVSrwkz/SY/e+bIUnI
izjswff9WT58qhNnSO6YZ2hQAb0xO/Tv0F9HaTMvI18dvzWm+NpsNb1uKz8aE8ed1iRuRCFzeD3r
E5H0JMbRAuVq7ke0b9eZRn/OT/EEN0Ns43+AmCpEFPD4tnZN6pcs1/A+V57utwG8+P1dDcunXWqZ
hN+HErXHP6VdKXzMh02FluSkAXhOkGJD2OLyu5MIjs8ssQoFS50xbkaNXhX/zGGDOCimlH360y+m
92F8SfjjZipuVgkLfWToy7uBBbpWPMkDi2W05tWBaUlJ3JvASqI9z8lzVvyeWDDeL1CVD3UYlnRV
BLuJsCl5R9UK9otyEVMGRD9NmQHuI0wonbajbSkk4Pd1MlT8Vm8iyc1zi+BP57Q7mpp9IKreGenz
hXrqZnqYXyup5EUder7QjETJqJQYKnH5LxTuFe7yBBdCb6UD4i401k149a0orobVxLQy81DKhBUX
o1j4zLeuklx2UKvdTMo0Z5NdsZWznLNWbE7UznCvJBziQz+9ZuHosAkeo6o/Rhxj0hEqa9/MTw2C
Zgdj/4cz0XZjcinXfmFSL+4DlExkC7aAHgPuxvnq84bRC60+WGsJFSw5FIBKC4XF0UAzSUx8gwUL
YS7uhfBj7DGZtkqp0HTUVtk18bE5y80ZErPMe9dW5gdaZHMvSswi1FuKn6VGA213onxEtY9Y+Mqf
AhVRrWANUDyDof7fGuZvEhtohrWuSq5U6nwA86QKtKxkAP629ziea2gWZ91SWL2qIbiEyQ3K+kda
e6xEBNQOOv57m/o9S/MdklVXlZe9gNPFH2JWCj1t6FroMeXaawAQKJY/eRt/oM2rVXRb0noikt8p
RGqiyhfQtaV9ZPQA5ZG39785hwZun9ukeD0Iq2Cbe4VBxw2Ofc5mSEeHvG+dxxgWJv3cquqCgt4+
66S9hw4rVhi/+wKgu0FzjXx4xa/Lp26AQjBmQXnKL2wHzndUp15c6SsQfjxE1M8br9sKjSZmo7oV
1jVW9uanX/BOZJSa0mMUkyzG2ffDYm6h4078P7qBMx9UdtmHVLc2VCjrmHMaSWHu6UWNkK3TKIX6
Oz6fwHfIqyGegQ3Xixq1iPlmlSENj3Zv1M6S7qtrimP6gPaNNb6u+IVia9frdIJbTYadMSALu1+L
rhMUi1TFifsMEzaJ7Rx/aWl1GfkIEZtwyyajVbXTMwDfiuRNDJrd1CICn9tWeI8grTWdDj/F1qZb
k0qlMZjlKzzoEh7me0yEc2D7tk73l91W5nozR4CQJSOWd5wECZevKONGwTxHPmjh9pxgz4FdbjDt
JfxgahlVvxgTK7RIKmpbmrEU+YZOGuF++3JTuujIqv3YM7OqJn2sflYfPsaSihJ9LSSj8hKCs6Eb
CFlQz4sYBBCv8m2qhjP3ZoKSM6RKWL5ZATv2F9kS7VLuGsHW8LflDLCdVHSl9aQmZP/76YQAJqLl
E4cQ9/JxK777cnbLdNmIT7F+RVSbLqsjkyz8tt6IDQZv51oO2DRrASe2dCPEcMil8QGaLGQvbahW
+qbOEgehguiXxb8HIrK4rulBU9L0kwt077wn4/4PiwaOdtrkRGBhbdEyXcR+E7BSuvcAo0jUb1V1
+/TD3cLyDgfTuaFuw5OSXLT1CKPBBOpz3G1nkc66836gNFxLR/7MWlJd/p4fl1FSXQn9aA6msKsT
09BvPFBHWhifY7Dd9MXEV+fW6OeFOLd5oL8acO+sQPchjtQRTh1TprhojB8aPq9LgddF/XYmqfQ0
rJTCplfLnF9gaT3OTLobGJ/JPypXd6+6tw0CTkPfS4n+K8nfdpx65/R46oR3Y/9hLXM9OdCdT2cm
xOUh46Q1T34lNMZA2F1JDeqSvVAyPJJTa8803ut0iKtDVMtvaOalSn/d6vjZ3xHmm8Y/D+UC4BNr
kOJFefUlg4pILb1cLKnj9aI75xKjOP08KV0hBqMFT2G3dnqjFC9LEr0oaBkxYZ7l/j9uzX3WH0g0
RwYN4rD5GT5uPL8KfmR6YwmUI4iL7xCmoRjdabczYyhS45LcOvvnmMfXyOK6r1Hn4q57PHxshknI
6GfVPNZ/GPz/pIMaklAqNqA972atEBvPrSwOXLzPn7cZCE46bI9I5rxWd0y2ove9sogy7dg0lA33
A8E6WN8EzE0AR/NnL8NwEsERP8hR3NAVcwcvwghnyi9E+joVaXW/C+hJl88JOBRar77puy4u2ndi
DSlNurqEMkZlpcncwjmuifOMFL5OHZGwVi0eECvtkLrTRwl53MmsolQoqQ6r6xCJ03njvlSz9HkT
3E2q1C/bQabYJKVI08eHBkShIa2io5EUXB9918r5KHxC0YVyI9Xb/z3ups1UD0X2YtLkrZfi5Xvr
499L0C2uSNo20Pdq39ZXTw52IWIHvm4U5D/9w9V6pO2SiZE2gS12ZImpxABVVScpuWagV5/oCutk
SV3TkqlDYsYaPjkQxYfOqXMD61cnI/P9atpUIGHxBry5PyCKii/v0oOwTf+M5Qt3vKsat8nOnSkx
LB+trXSdx8Od3a59Ptr58WMxK0bxDNlfhZ/KOY5pl0kFiXlZvLareUl/7oYk+fv0HUlpZrFnzfuQ
qurKKsxRCGrk5JdUu1T2E2R7FGrFwTvtwVVhtQPqWdo35y4eeU/4x+PHgT06XBAJHvb9iWvpYyQQ
txbMrvh+YuGWtcK7g40zc7ccf2nSKgCoF5/R239EwWF6IkBeQ8A8TFT5AcXxRmFRdTnEfKogxTqd
YbXFUzXWeIDDSUCxYwGg1Hdu5wXCqTsL3dWcD/2RzG/WFgt4pXALQlpTZIXoBrRvegyiSxEaT9t6
FGLvQoKEsgG2ANP0QUZGHx3QSPOZw8SAij4fRwFdwL5/g3rzPs4xZpCXxYPA8XnfV6rbTGH7PMpS
rUG9PxOJ2BQmFqCsejKj3XzD/yOc7kLcAVSBqnP3+x4Nec1mk43C9WYIop195QQcEHr19Zi0flAT
TYrI7buF1XoezKYVJX+pQU7YL+kckBWSaYeabvJSq5HVaRlFLQCOPgjdyVJdb8OcznYknrQ99sBx
WmWJiSJ3wshqqBZpmfK3dRWtYeuoC2vNzERnGvxAZ4XUyS254C1Mw9b7gmfTKSJiZL7QWq78R5zT
7nTsKjFs3gxEr0nqSVUD4A+u448U0z1L1puf++JikLzY0uM8IOIRhqtkr9T2lLVdpYgyDSs8G8jC
e9YB33jD+bg72v0zd0xzOmzi8HQlcWGDTYLz2dsXVp+Y/8i3Zb3CSOOis1V93J8g4G0bNTqqXWtA
TnkamuJhawCXnqY1y6NNfpqq7YI7orYKlzbDrgfMh8ZbF9Woj0UGDNsZBIGgj46QunHwHvLVJjSc
2L6SLycUZSIK/ZGkeWHx7ixKWpMVGPATtQbyiALNrTFQaoc0G/8BIhz89Sbo/XJz+5Cv8RVo02ND
ik1adpFcB3nvaH99pKzDQ6g0zr9EW3XZGqOmO6ZcPQlbPw+doFpwfWMG9B6F/XuAdvTN5G7rHRNj
KXnw0uHCKSArqSNCVMnd6ZwEsLHBabNzVh31KjUtm6ugb07OPv4GW2kc88uIVsucOznR8Pw3Qn1W
YHmUmM7WBPim4+nugon1ZMKOKQvP8qpjftl5dA9xsW+cKwQC8c4Gw3f192wOAOOldzGFRy2cKNRl
tX1kxyiYJR8i6paV6StYlviPsEk07kYNe2OYHwsaCef+MholtD2pyWro9YYHnVsl4t1+hxOT0ll6
1cxN9qbRemSlPYZVATtXwQ68BGuy+yJPTowREuHHSpAmFSvfKrxmFE81/s7Vca8BYHE0jge+VMfT
i07t7lRkRVmX06Lih/jJpiTJVZks5dLgvi4KxsY9fiUhTExvFe36IwqDyUkuHOetqUKSto0nzG+j
BhtXwFpPnVA0GvdRFmgDsQQFZgAe/5CBXMC8NQ7Gs+12/5pvCWU1tJ+0eX/NJbA5y0m0C148X6Zm
3J1Bjs3IwY+UKxNi1ulOAYlIcy5HIxS7ZFGctySaAAHex0HqxT2ghMQ4PfAoHML3aTxA9PXFjAhc
CQ8JVPfktOumdiUArMAf2fLWiBY7nGQ0AHl/jgQ0AZcqqI29rumsXlKGXFeod3DVNmx7EjXj5zLj
JmLAP0D6VZ/TJEFJx89Kz3otMGMJhwYGtkPvMPY+4lZtgfMuXGbfVx6IWJid+oJtrPQRYrovPQFX
ulgj8V9XeUv+edRG51reg6OIgw1g68Q0n5aCUGjYQwxLcJrS07nmgZM/mi8xH8/rY0uLolM6CHKX
nGOAyz5Zojb2EM6imyNTAHxtuyGvz54/FgbW2cKFEHWYZMkFFkivCl1+X/oLKrWzBedkSOb6lADO
d7DRgvFvVfnu+C0pPgQLdRAy3mHYXldcb3gqWImFZPqSHggJ0RMRYo245IJOrdLTpFHWY72JmKhl
oJgDk45xeHq8KHptwgFmU0AE4nZO6Kppm+edw/R8+gmVYzGtJUTDVba/ZmdH43r80wYSW/wTgb+K
a76P9ABDdbrx9kYGjDYboSnzzmyl/4L/4Gu8+dMV9yie+4uLO+igHo8Hkm5siR+lEsF8alWvKO/f
PGA5Ci9qhv/uta1ha8rLWtJcIibSxjqPTglwta5J1ZPAd682AXzZ2X3Yb1fPxJlKO7I6BHszanH2
dR9spd7Z2OO5X7R380/E30Ws1X6pAPWfWFp0NkKs71hQOhYCtLD2DbuUg8OGuzNh2cXEShu303Tu
8sQ9lIfEW/cIgzSzX/pT09Q3Oa0Kj4EarEY2L+qkBITnuxnO+kEL+WvzTrHPPzS4ZEtHksIseUfk
6UCN51runT8BQUIItN1BVkGf1tZGOYdWNeIi8Pclax7BfqdY9tzG1iQRhIky/ucZEZP+PGVSSA/b
tzWusmt+K21DeXD3iSw0PEfDfS87BHVk8q660e1rOkJ8vsT22MuQxIGAew0PjrAAfy5ksZgLBBZZ
9iqaAuKMAHhpCKUAnjoiiGPvnUXkLyNXliUlPg1i2bitcdU5VxI/IOkEWbJo4/zK9e/fuiM61D9A
lcFzW+pE+OlR6Xqbz2xP6wm/fYwTeub5NdMzlmx97mpew9BMnnQQJcIwPNOS6pT+DiDxX5ngF8qt
66A57ZJOjqRQC2OWdGi/Bt8GPhLHuQo2vQnDH4Q6ZGFK7EEcUm4wWo1f0/TRzOqxc8F8a+Ly+tCO
rWvEPaORKbaKQL3IvJpC6+P9Vl/ZWi7Ok9YTGfWRPOnoCrKdShzkA0KtfIiW+J1Izo1PYicTJThG
7xvSdyKdRtr5PsuKgSxe/v0ZM6LIdVP8ajpppohsHVsX76TV022IjTmVEvtQaJyfMhPDBBvA6+pd
GfDzrACkTbIG2qOkSGfKmundQhuyGbNF73hAusm2ULp1X/BXcJP6ZLuthncE/KAYsNlp8s8SuD2a
qSxHge9kEmfJ0NKs0n5pgyTDr1KnQeduchG+syI3VWne3F1mIuX/qn+yhL9xTt7DbkCUxt7Rj7aR
vNu7x3CS9SOeB5XMO19laP9GkwDERyfaEPS95pbErsyaeBYmk3zUvGYjC0xrtYSuFEOjkN1OcEVa
0UNkTw53T4SSH38UoHF5Tu2xQ3pY686rGIo1TPFxa4qtnY8hok4JbHb1uxWp16Jt4eiWJRmh3Peq
kU6h72o27nXDjze7DHVhazrx16Ad+L69q3y55KYgmJIWoEcF994iTviVihdx+wlF1UWHVOQCfUT+
OFHEXH307LYcCeWQL3Fulv7kcH6T/9+/4552IHSAvAc1MrufH1+OF4QagDEm/ATaif9SH1OSOTDu
un4kz7N9+DtqdVzr8E1njJSU4EupeCqb9pOmQSfAOrvIkr/37qiytbMPjrOuNyM2ibmiTbLGCErM
mbhWbPC21cuh22q3VcN66U8KoykVhq8wwOSiwL9h+Xd8QU4faEpeJyfBcWHzJwFnH9zZ4CsZrmoR
rN8D08qX+7jleV8NbgK4+m8P8VcUZCsyWNTi4ekDL8r1yxS8BGTgWN81kUyNG8sRWqXlAYW2hlG2
Hr/u7uip9pQURN0fOpQ29gGjMJD9fduPU3eoJJLB1cubKd9+zB7zbUVzc8c7AIqfbQ7JFTUVHQIs
pLv4w7JndwERfZL/cM5WfKBCjEx1gLiTlTatdPi5dHn3oxtJ+ciOQWzyHTuLZEU9rkVE9EO78FwE
nclmQS+VJRucy7JFH16CH/NkAorbiZx+N7N12njbtd2JKveKglp00uyMHUIzosrXjkoRVBXTN2a5
f4vHarTueuvxkuMetVw2Fsyw9m9OMyvh0pacKM35TTdsnYElBNe1HHvlzLwDksHeLiByW7zzBBC1
k3bwIFcDbtwVq8qt25MaaPgPEi6kShAQjCJUtnTGcu7SZscBD0EbPqV0FIksFk+y7U7kgaX0bjjh
JwHVme3fp9911vCJj60sYYpnyXU6YnSeQFi5++/ElWoLmy8lpVkeYqGA44nxgPptEz3SKUY3k0oA
vxU3VGI16wM5GhjudTREyuoTGV9AuEEl/oSK2QxNt6BbKEyDo4wl/H/tyETPIMvx+99VzvVxjCSZ
ux3CVYPhoRF3uKeQSN2LBzC7rNkpxfzZUIJKw/SFKFg63pf70+JbrBGkHZ2fhXZ92VukRB1VMHW5
tvh8LUKM5vvjTYTzG5pOisRfhSh+zr4G+DVVIT4qVKbsX9WzIIB6brEwVbv4BDgr8iBdGFrEcRDT
2WSWPcbffyh14LgzOdhu+0+Nnt34eqH8qA8pOGdeOUolRpzK5H3AR/TCDdV6wY6e6UQFaGPYYC0e
wYsruAZnQJtusT21tVagHZut9Ff6WCKT0mmWjy9ki8MGXd9LMKIjikr1OkeTtWa1seBDtkdJkn8F
BBTn06Db8+rPrc30rfOggWQZdfU1ax1juhRtPJWEUIoI+3BoLNvFEiWdhOeiWhSKm34XkavKpLRT
872SydGpk08npckA36J3CLITb3BIlinVX3msRp6cmtVVynQ0EuLZgorH2vBGqQno/A5dOGvkWCRy
0CgXPQEKt6XWAegEp0kf7VAXREjBryqVOzKr5RauNTpIcgrZUBFEatwk+T9wX7FA6eeXq1Ftrc5E
hGmRJvYRoP56IQU1C1cm6+udeDQz1COhvVX0L71bYuYXpRDnH+0iD1RzKO+KGwdBatV/n8muZhpQ
9AFhtjdkhELz9pP1zDM+M/2Q8M3fjvMkwIPKVW40yUoxA/G908xKk0XaDqsFA9Bw4bHwnjn+ikT7
zhkSF1tPTTJDqUFz5Rxo6XO8vUhPMN9ofLJHVxoxTIO1UQ6lY2PBHdigy/S94EeyR48KDTXyDOGX
cYVgSsX4yA/jGd8UqqwR09odGzqcOym5uT66jL4aE0amBar2lbZhNpzKG3d9DL/fU/OyLzzNg6Ac
j45IWzLi4s/UQ8ml8Vw0+k5ewj4TtQ4m2/NWLNL5ac7h3oWargfdgLJSUi/bRqPax47K9DzKT1iT
utIiRIZA1Wk6TrRdnoyoS9XUPBX/DVl7VSmB9gYJDKNdRjS8pxvEw7AhldB4r0AoceXndJ821o0Y
Cp8ubAp+3WRkkHgpFsK0BBxA7Smkhk1gpMpY3Duxq4p+U5x++2HtwYaiKqYRflVBPvlpnHAFQKF/
DUgEz1U5CNOf1RupXTO/61/F0gFEqKt9QDMXnSdO8jmCqxxf9sF297UDcTPV4xzLalfIunOKNQ7T
V9C77O993vuc5Uo2btofDMeTZOOedZA+ZOpC0yu+1SBDN376ZOdaqW6Dzm8eP469WG650X4FinsZ
q2f0p9SFNUVbwFzdmAJPAxXiz6xVMPc+6DZiaGZFpt5vGz4LCCDT6IGAo6Wnw4XUAgK4EOSVZ/B5
47PTut9/FKWYo1n85IQ6a2cZFMfrJZafN3YDTTTx0DkTRBVtVdZU8OMsoW+QJOCMQxAf1c5rP1SE
xAmnqZb8zv7ZxVcueBW0YOKjZf4141ZWVAnepoosYZo5Cj26K8UqqI4Ln6R+FHb9tK0yADjpvW2E
00r2SwlGs7oiODTELjrR9cEYT0VRb+OQyzEvos0LAub/HRARV2fdirYIyYhwUH1fuVG1jq5pmuIr
tNFKO7ind8aYiKzJjZF1nBJWw2+4j4UoxBHrGTkdISn7oUddHhc7GErO93xqz318EdFrOJkIAMdI
+tMKxYstp1yxifs0j44xMztVaMFDTzcDh5sXDTgZuWWRYHgIrEeFo40P8tNElCNlg+5AOt+71YCV
2tISEVFm79StF4mQrMHvKHL4vQdRioQR1oCcIcMX2vDF2zPDPkY0ZeVdNkMzKop/tUgeN+P+FH23
aN4TrYMdjaK7SqR45vWpgnWe0C3LCTHT39fSeUL2WDpN8FqxwtcB6+4e7+2AFzFhB2MaaQrT1qTw
RZjEod2oUhVcCwv8qandh0S0ZEWxFiYLiKlerzMVBvPP/NQs5Iowke8LEZ/braAbnNaq+PP1YATh
tz9x7rKE0zxmqfamK44vFKZgohu8ArQsLPJEb3sdmbJYR8gG49Ix23BVx0OGQrmoOeOuot1MqLga
io+qoMIVaykRFSECmdLjeR8TrFu8wouYW9FMerO8Xc3QiqDQmcdvUU20ZoP8h7CC+KF2yNXCzcc4
kVx00uWCNMy6P/CTUiQ1U/JmSEpwn++/iafSKYJOS1UYiZn1z7J2SmE+Dy63HvGfeaQL6EQuzYgK
qPzc4JO6eRAigWp265fkk0tJNKxSIg6PsG1/NDp3XP+qUAd2TttA5+MUJvA2njSO6fji14E/mqje
kzu19eCvNesTL39cV4z1gzsrDPut8oQFWOhHiqOfbXfDhSpnebTKTpUnA3KpbMteqMI3agZW6xcE
NF9KoFuQqoHwl4pFj3nYkqHE2JQE3L4Ywt4BBzya1+klGibSuIEDDWPzscDBoEFpXQoaHo/lIaCa
oavyrpWUKthpzaR+f3m4RihcYA0c60JFYlFBXNOuKLKPSIyidPZliwdFc3+Ja6lY4MIMxjDRpshe
1INxIGWFW2AVYBSsI+bJkzVAs4U6RSFCCoUpGa/wfXtxX1EKB4G2nS1B6pz6fkW/npau2YYwp9Ux
SlzFLSK0lnB3V/rkvDTtV+kbj1oyMKJYhA147AWb9+KPQF9r3TOI3hiylhYcf2dW3Xy6Z0lakLkE
h0TwcHOrFigtqe6el2DiaTGr3In6DfPT+amdeGVYu4NOd065cyK+lToj/n+ZtKVzoBMmsTwRHrcJ
7o1DrZueE+XHsXpuetLbtX0v54Za2s/bcc0M1ar0zWzdrDgv7jN7Xe8M2Ujf3L+lbBOD7B9nVDTD
rfz7xGBPcWhHtIJbYYCJQ6Pvw14I6zbdAyBtF5tNUCWXeL890A933KiLYKrNcxQkcrhjCEokZGGQ
k4Q9WoWl6EpGQB/u0c40lotxPKf0WXPtmKb3GF3ZU0T2/CLh/mLufiirz7ILmYBeemnXNKRRLk/m
jfIl86j6n4A4ib4JbagKECDVL1VSzKa5k7QicZr69AFiOYgP6e+gxLyXKycgTQCE3riOgX+5E1/a
tzvzALt/QdW5+iWv7bnXJ/kuGZUUoMNZvCLKkJzCZoKxZpb0lS5jnU4oeizt4WG1h0Gd4WDOYCN1
o1CrdM0to7MK7NcckbE5t5hzCRqmZ3kKgdGgO67dYf2btA9OGucC6fyk/UDkTyBAeXI+rGOBaQuj
X7aBjmRiTgk7bj6djH5IaixkJL5dD5qA3lNwNU3cgPqWYkniyJI6WeVB7aPV6qY0mVjyj0iyNQXb
tVFHYaZqjFSrJUeHlDwf/nBhCvlBeR7XK/Yj7FmGMTBDwnOoFL6KSnSHGYSGy28QO7o8gNZrb0GO
AhD6vOmp6PcdnEMnimIqVt5YeKiiOWRkB02I2B6cZG5nhFeKXjgXHXAsgTqf8b9QvJiKw5GuEVDe
HYkUHkFkoBWmU7hSQEYRD+Ge6QxgwJoEHRTh185+BFU56Ba+/lFG24cLkMaDrMvDMCj5UxcHXr6+
gV85eHDvSDFaaZxWgr+Ut9nvNxNSGe/slPhuQf2yTAZO2YNIfzuWmAezrAuHylZnAJsapR+XUCsS
zwt1emuTtVRxmYFq6qg7x5KN2dnHNgLAr9NtdiBlJ+lFepfQxAUX+Ur7W7yObINc9fKf1oEJjk41
jsVxz9aOpcOux522lyjgSZXFviXAfWolQbxLPe/aI5YDVqLWBdYQew/Y/Omb6PqxVTua2ckVb4yd
XgSjBsdCE9td5nDFst3g2pSUd+VN609OXZIyxUg4Fxg5pyFUJcbILRxl1t9byzQb7f1s4ayVqXu7
g2v5RU6h5REJwGtYaW8KAb7o648FRceSHvK3LN2VqBe1go28/ECdTeahRR0JPqKu2tpTKcBN/Ybp
3sHmGpw8e6tkuwnWsNtpEGpkh6pvyazTbIRC4CWrrobMne1gu4KZcKKzyq8HYXzscyTCHdYtPN5p
K7XBKU1XjofTQ/iL/AdCIf0iVcyl1Nq2ZYBRsZKePp1XmfP0KLhY4b7t8bz8XbKj3uz60zU7v+5z
a+t6bPLLlwP+2Sj/szkY2mYrZPNNcOLtHLRRTJ+XXJe9AEFPB44ogOgBuRJ/1zzMXGmOUmty1bly
ZchjTjYIXDx+/N8FUlpFUD3m9Imo/AzRzGJuw0jz7Cqs4O2Wf/npc+aHJ0Gjn95MHp/whEB928vE
dKHJzsNqWT671ECyZux5LPK05RzSHS+VtKoIDJSU1WEaKx9vRikXhk6bvO0Lcdy++6pZdkj3LXqP
tXOb8ImlvkW9x8hU92MEjQ8oPXN0qnDvE8SsSf9164XrX3zY+G2pd/KcrclYNpv7sCwQdE+ZQ+KW
D4ao55OwtwpJQrWqItPhRotpQ581MF2tPYg212qnmSSFh1hPBKZmvVU56fSO4sORZDiAJsXJAgYj
SF2iRpaSxouY7JpvkScZr+nB6Sl0pD3rIdJIVtL76y1qZLynuFq2iVBJQ/38BxF42FB08vdMDUS0
Fy4h/Dj4YqVL79cRWCo3WXIDEeDKaPJMsppijG6AWtgIwLWcJSj5cixKFa2DmSiwcSIMifm8tVYx
kXGnb0EX+id63KZQatCwOg7sS0LAeE5K/h8vClv102qQsb0q54aiNBCrkWpuLvjzdeWRQJ/CIe4l
Yr0TiU2TMxn2NBgxg+7OSJsuOSqmih3P3G1uLvHDa0tv1jNAgEeMfXzr1PbxldWGin2WSjb4gagy
F/SmWWLmVtKcmR9Di0+DedCetLPGEDqTjstW5NdMOFHtLmybWjU+wJM9Hlx7oVlTljAEFMLgbxe4
sqMSpKlPM15dUnJPOwKksv9digmOJMWRQC32Lgs3frV9BkF6dMAIh3QimRait5PILf1AEbqz5hij
CQnyuyt431RfRL8DwDQHNSo1uWr/bRboAZfqIofJiP6mYo8QnKhQJlzrXSO/fHZTlk1G9nPyBPLK
CVN/JGuxHy8y6tDbi71Aqu8WyVwzpUoHMnJ6QwinVenOKcHDXMft5z59AmWBK+whrfV41yCXM/py
hY3or4vyTzBi1KXI3rl8rbTIOkB4LQnVC7U4hSgATnWNaVbICxx33mvCbwQyDVq6GLovjMRPWHo8
UNZoG4PWOFfYYKggHAbWQGx3DDXASohegbPbrRDP3AiGyd1haV3zmzBYVlC3UGuc6lAIFM9KTmGH
yY0Rrw5h0wnjKvm61cPGR5+JAFzbPpmp/v3XmWz/NOAV3SjybjBUAKNxR+K/mMQQgE87L3Lo0oT2
1UXXE8RsHWuEFL5qMBzhB691rHqsOCW985TFMhk1XrJHHZ8q9OqfAHV2rV3dTkuWfSznHOpoTiiU
korFqu2jpai84PCp47+HDbR/D0eXfKJevOPUuE6RnCSKE4Mdq6bd1uQ0euY1gejF1vGILcBCmhjW
6uPmZciLzNMFAsYwQgcpD7atem6+1DlO1tZzOI/SNpYkUZUs854xHSw1EyB62yjijwb72oproDTB
mVw/20IjHdtAvigxC+kq5VAx8kVyimV/O8EJWTJc10Y/kGHu8d3v9A5H1BKqiaFebqtlWqVGjFJp
oms3Mvu0rQ9VRljLQT1OdCyg+wTeGW9mrv1ZSJYez+4EngG1/Fx6a8nlnecFlwTODWNUAosJjqx0
5MM3xa34cV7ypzzgVyjL+ofD+DmcDeLdZSlXzKKf3Iq9pV23LiB9Kyn2qaC0xkQY0J8s4XRYkDYv
Msb7W7NoGHkUDkKttHSHojpMnjaotYamvQXwEkxywTDZoX9SyIBMTQD9PO0o6jsk4BDyM+6Nnv+m
inzQxi7hK5sxVVenuDK7V2TYdBR6jj224azZ2k8sKwcV7pK576Q+VUQ8QKowMmkjeqDL/ifbexZy
mkqu9vNtmZCVIWn8yxXlmTpOpAQV8Y/cvBVa6+iyVK7/ciTKHiJxiwHSF4d/XxHPiT31IbTD3VC1
Msc9UlfZU9bWkZxOun025dsIFyFBofXK70tq+pKi8QfejEQqoHpqMPoohzFWofR1hHIbMK80Fxvt
uH4VHchnuXiplTItpPU1UezDdWCdB7cQ/QE1yfuKcikFxAIduMItGTo0SKY/8kHs3x0mlSsbf3eX
vNXETs5x3vrFoHHmWoWDSEoGHehI5fckGlGQq+8brH9BdLhhKf8Hj4yXF4S46atS9jkWSWsnkioy
yVAgMUdKZo/+Xs1NhNjbwixS75vfU39oWJn2EIsLUna4GZ2m/A+7aifzYQJIjwnmKQ8xOTUh7Twu
FFsPV4ZFLfGVytrN4ADSzGSGhv5oksnGo/W9gpwvL/ICxOl7S1n+Q0ns+g0qUXIwEZRvOiK9oZJj
sneJ50FFxkesjzl7KruddnBVmANSpxsEJsfaSfpISUJ8sU2RlaygM5ZXwf9Zs/vYWfvgjRgf9n+O
gqHxsBGI6wafOCE9zqvPO533mX5scqUddhKPp8/HugPZxJlob3HUuTdBRFAFpC71vdfDU8aRdQCR
9r8/l+4W1XtpKENDt/aGhy+RC3rKEchl9rXCN0RCol/f+hKr4ilfnSEGYKdU4A7kHnD0ofDsg5Ps
vCJ1kCN/CBnUABDa+TpzAYe1n7cIEy3CBDMDTx7iXi2l7CV1untlahNdHkT5CoDuk4UW7vRWEW8G
/kpTtzWU5m9dsjlnjqLCmsoDM5JAv9C9dtBMIQcs0dDjQgzmr/l0jHV8ydR+KCZdIcsnt9gcVr2L
IhqQktg47/PBRwLdhhwSQpnV8OlbElqcPL2jtKVz6+BHKUDaScumWJPuFl56OJc1EJaOZs1kbhwp
K5l8Htnr4IoZwro7nAv+vevy5IBiUJtc3hq6P5zj20IIfLtw5nZ1onwLWNCUV+yEdRFyjh+YS5zo
1EHlRuCs2+K++c6LRqoV9DhcQ091inHE44O+LATjvPlYhIiffeAqIlQbH5P1LuczxMnjtnIW9NNW
PscuvcNqfk6MJYlWke6AHU682WkBqSF5IBqE4cVrnmqYGFDVonUnPOAOCLjhYfVntzHLg2OB6Af6
O6jnhaScc+u9rdoTlT98KlitAAJuO0K1Lh1bGZ8r8JWK5LubPVf77WPrY4wzPoNJSVbyDhXS598X
7pfR1boQT6bmhknZYkfXFsA+Mba3Uad7lz9L19lMPoBmAol0HNbHL/jX9jixOTgwTqZjY4JkZXXA
2uVyVRYFlbLSf7MoNVaE8fDQdpa+t/UBFJIeU9GziZzxQnlUqACb4bXCG6UCITcgJ1tq6rTK6UBd
Cm7/7twjRg22jUPY5n6W2h32T64tQ7DFJZh/Dyrm8SMCGjnoc8l0pkcHfZTUXH6B5A40P7hD2ROp
EvH9A4hANP2wXgCf0+S5+cs+SBwy1TY7i/UtO9PjVWZWzLvIsF2xj+k+fBafzsMrPWnRaC7Yo01J
/6ji0Ee4gN8MxAq7BsjfeFK4Fgq8l9m8h3R+KXpZO2qozY6hLRNYP31Qxp9agCvL+P85NKm/iCKc
fRGlxrvFX+egwXvsQib/trmUniaV7/U6tWDixJ+spJnsPJIY9fXrRVOtIGWZuV/Z9e2lShg+IgTw
B19shhZSrbW4t4s3Zz9HH6lxg3G/9cndU+DJvL2MxkTfzKFJudPLarYZ1yDDZt52zvtn0e33SQZI
7lpEKqp4NgpVcbvYqNcDkI200mDHcfQ7fnvfrub0AT8mJygSxD12rQWZ+HsM2cRZ/FYgmVAyLT+U
sQk7SCeFewpNVFsTVwRjP0yHXyx2ezw3hThL5gcY2IZV4F0UjKiU8VVkEAIlGLDz/Mk/OKloJRwB
II40Xoz19YNX4NQkvyLtf9TdLdUGR8g6A/LAdwLjAPq2pCJVm3BqSEmafW+hGQlKcP2KWzclGH2S
K17yajV2BYzNDUEHFE1pS7tmALEny5mrtqCfXQ8eyl9XdVKCC7ipM2nlzw7fg6WKjgfJx5FFRMRd
lhd4GzsD1AXWvHtAOAt4mfLNrJc5sYlB6d4M+mL3XsHE/a34aGedyOGdCC2GTD2EHFQVK5pE6K1O
T4fPlJU38l9vxh4H7MZRb5jdw9igF/zcGTFYbf08+ewMdwRqTVIylKYo6kVKJHm9XDBeWoR6gTc9
h0O93fxG0LXwGmxwG11vVw/v8qdYIuRHcoZq2HF1UFQsAq0XnufzqH6l6voDwPYBFtLTMIPMY3bu
wrQQcoDO1XMoYROGKPM9OLk8A2bnnscchQTYg74FO8zlkU4EvcSVXzrFaT/DOOKBdXxHynRC3+8O
/ticZ5DkRnmcmfbzdlaQEA+6nPwa4j2Soe2cqzA9//zfX5QBYiNadDltZHa6mKMqFNRGmD17RiMG
B17XZFJZKOvLqFJWo0vyAHN3Q1TN+LKuB1NzR0A8ZlSZY9P0QnMXmH69e3SmWhhGCKi3+uwX3fIs
qjFYTR3AhRvNcertIfMug3V3vAnIWqV5mx0zZFtzdpSMzVGLBRR9qJjEuWe0HAim80XCjaILrlmP
vStIv80SK+5hlYX4tdQ5ZBo3kf5lDyMtD+opO995LSr7tojdHmJ5Xh9JNVh3x9oGqSnRd9f5izCm
HF4nuWCVpZ9MfSXKibmqKfUBYaGYcTbkZHb/2+OHpN1BlUbhhNCl0McVeRSuJBBFImglC0oZE5ra
enITWJtSirOyiXnJyFUyezx1hqpgW0z5APF8u578S0Hzff67G/mcT1cy/WGFC8zApJQ44kMX+TkN
kjJgsXN4/8QVaJE9RWcdWyVOJmrXcqb5OOXRCuBe6+FVYWXDf6LHl2Pxg7w/U6jMZpMIlbbBsh7t
CUHF09u7k4ND2Z+OGEViVGcG//ORIKJ6pyKvGtieEG6Z2bOHdubesVSuMj5ME9Vq06nJh8nFaQ4J
+k5qSikvDYZTRegEUJ2PqiPVubcF70qiJz8j71Zah2/WounmrkuRULZw/2PeY/DNIiTTt6sGIZUN
gc4aiFWJditvbQSm8wVfKYkWSPPlHZLljNzfeSXkt3iOJodiJQmNbaMm3Xi9pJukoPdNHXCd99p1
H0xmnsNVm9In0FLSKmdSzPclKK3oGamI0oPxDji0nW0aL4kY85XrYDuhXBRmD4pmag08hveroZBy
nQQEdBEcFCAYXNXHF9Rit/TMP2mQqZ+LDKe2n/8oQCztyOh9o3tcJJK+Sh3k2V3S9JZsG4KpZtHj
SX8H3TJJpa88GhTYkNupn2A145zSMW1IHjWypv+Zjrfct3x+A257pmj6NtZ0kdVrw2yUQB2ot2ay
oTWmb0nH7n1vsKIwOSQdK4vlArG/r8rqdPP5pGkxMS5YrtnuBCC4XDu4TxmEBxYz6SJulydoiCP8
TV5IPpmAjrQ4VRrOOot4CAHjnblYrSkloQlIf/rKH8voWz84V8W5OSYeWZpXPM0v0p6CE9O2LJLU
uX5pVf36KzOwahY+tf/NnGYPZMK+S/WvRVTDG8We4fGVd64TqZdmA2SGq71puXMIgwS2wshhckhD
MXbp1XPHz8t4JJS5fi+ult5aIjb+4BtE5TsUSzrLGXXaDtmRKZk/PC8OTWLOrGZZBsnH6sGVgNfN
jjAnQcS+KVpzgvpj1mXieISGU0+qjVNXttuYriS+GIWjh58Ylh13/SoH34FV9o6WnuiBTAoTkqQo
euAsTSkzP119dK+VtUcRE+jyo13SiQjto6cZ+x36oqe+YOROnZLdxKpvPCZhPIZuvYfZXWdQJDQP
OtrAIUQyRtxbjfDH0+JX07+wPVKciBqtwd5fL9TsPxQJX57+QbkWzfT75t/Wg9U6DURmb4o0XOSJ
rucbjD63RHIsE2I1UzB+YjeT4TnO/ZcSlRwKvs3xmt6RZ7TQ5GJCCv4q4PeDl7Wpyx56AsFVcqI5
q8fwnrEKHCUbrzW3v6DNCB+4oC6yH3RzDEBjUNmPi+1yxpS/PU3zv+KXtihPd8sWb6mJKfBFRrSm
+Epf4dAI1CxKseb6/DMZaytz51/MJZ4sa5ai9s8TRQ37K3u9sF6wUxru/xNmbnEWsMeFZB+bJS4+
nnCvH2fRShU93bwYcVPStqjd2L69Wo0y/GePp3nTp7Pk6BZV5x3PoH7Y2ArjxpjiJSR8MkyVIMXV
be5oIrmRSQnjEdX7PO3BJV4e7TxOoK7Y+ZD9XoZQMOn7O/Xd+4PDL1ERsmia1bwuTlwfIFqVwDXy
LwRvRTmfK6ukdpRZ1L030QyFWqrwGXlqXPwSw1gdAeZf2BX8q4SADEtsa+gj2UdCDIh3u7KRflpB
wCNPZLw1FXb8wLR+6PpWAojL1vcNPUYDHocSphAkS8k3J+LBzUbKlo+/dgXNSUwwnstN8rFqdzjf
ix/59/8WBqx5s94qcY/5MzSTuMsaJvMB8JnLrn2ofVritDuiKKI1WF/WSr6ef3v2LvR9jtBqOi/x
dGjCEgsXxKXXtXk99nOSTf8BSMszPjVWEQmyzmHXvf1GfQveUjr22nD/lcOVG7Fnornuw2ddc17x
bkOrNLIR9RHMrQ4NzNOOqZL9RlsJ+I6LKWZkcoOygBQdgRAX3SBsucilUWB/TCby+g69Om1IKHN7
UKBZqzGX9Ta6F/xHxP9DnClkRXUd3jpdCsdiZtbvXPjURzMBHJZprAEJOUjtAq5IaqDas3LiOUiI
fFtqP33pxbaGpYI3zkR6o/W3OQqAA1mreDXNAe2C80t1nFIQYwEpaFKamYePY1PFGwKF4/9DBl60
lz4k3YdEq853Zk3JFjZ2/sY66QO+KvIR0TnA1W5m3JP15JaD0nd7XnmXCJN5s0O9Ux+/8hg5GDWP
+oVfbCXWrSlBEVA/eaTBifnlmQ3cd+pruPijarUDrCMbPIz3STZoJv+ZxTsJv1tMdHEKWk6vNzJU
Q4KgHR1b3HUvF4V7tdDHMAjDyq2/1YNFijv5VEXfOy4SWrkaQcK3cW0yF10SaviVX7hBRnTv1L2o
XZLn6ty9tlKT+/MKPKZFWGP7UoQ3OEW0htGu+jpiy2Tun3h3JuPzD1L3V5yx02Uvkg3a/9hU+2iz
vbbPDz2yQSFtn/EX8zFPr0Kl4w7+t5hPhft9+dOY3XL/FPQh5ciNE4QEnmOBeDKTx/dim7fjkdBv
XdbdxCSB338bdeid4d2BCPC3jqWOOKhuijA31TOsw4Ceu3dbyimyAAsu0Kt82wprBVMUI9rrX/k0
++N1tFKeGzB/9OetNhCaSZKxrOjIgtzS0oCoZe3ah/pG5hJJ+SjPk6aTETqUZ4AI5p3qLX0fjwG+
7Isqk7k1iItEIDgucp5OL9DDUc+QEnAi9LdpE6ka1gJFH4N4XNNDhS/uH8AK2q0Ry54EKSEqUeFZ
UbwPqD8KYooQHq+KYcIRvwFdHi9VRT2PLLouTKmziuxa+b3qQ/2yfsl/cn2GzElFxEzAzGLtMlCB
an4Z6/7owsv8TWanpoYB3xIRt2zWA6mM8LqpeqxTMTfYaKrs2GheX3p7HDOTulrpUCVpeP4K/TEL
mWvvdofSFH0EA4xMayi5S/f2lUdZAEBUVsqZQ4dN1i2iAxkLnKmfrsd3naWZbnqa/ABTn0uuL76T
n5DffisjuQEJt+negw4JrM9sMjvI3y4sYzku8FG/kc25hGT9JNh/MYgyKdnoVk4WzWpaYIHwHzJQ
I/MwwiiV+LK9FbJvStA80+Z2/K86NJ47gj6E6tY1ss918SWe9pTU7W97fIg3B7KYQgALkdA0ovJT
loRXpFCzTPHGiSxg5x4MqI5xHc5chqfVrQczBgQ6n2xOQbJbJrS3GMQgI6gmzSRurgUgdAjyxluN
kaBGp1ym8Q3TbbRA/ZufOv8gHW21oix9PDuWHDu7KAmCPyS0y+sv2BpYl4d7eE0fL8eJEdCImqeJ
nvR80Ovr0p0xoemS9ptifzpJmSQw+/PKCkf+L4V5dni1umT98Bo+ahk915jaZFHHNbNmK81xz0Le
PNDlNvqxZES5JRBeQWiMAVUm52zFqOBUYBAXQ4nqw844axMIja2wzVUTs8wYmgneb1BvCUp6Q7qa
yhZB2YydpC+yjDgf0YJHdao7jrlZef+r2lvrSR0zxh9W0hUZAKCFSMhOaJXa+y5yw4euj81AWqFx
oSHolCmERh5432TExAVnoGex66c1abQwoQl3mGfLcfjx8lH+tCiItujhTkgOTnGz/1srR/eTBLpP
suKac9BHB5WIWuxkduf+4V7qsUfLnWOy4aPgeIq4GqFrjGDxWcfuUX/2J4cbGotx+hxvUHnGTXfB
62Y+vAegchnoSrxrRIPtyqniGWRmWJTJ96fk4EJpGYOut2TQrCewScIvv7nc6VeXdiwGYsautNKA
5eO2jFnFcFzVIcCo8Qfbog3XQkoknCH42sIS2AiwoZGcXBNxuIaqYVwBODWj8bn1etJLgBfyEJ0p
hWEaRrGHkHtLva9hz4re4vLHITozfqXdbsFcn534qhklzW+6i/oxhS29mIABPa3x0yX5PHnL/hTr
nS5hZQsoMZcxLjx8MW2/erN6oi8162rXXwaIPPnUNmM6L6DCaMzTj36oxX6RCGDp+pp+ct3ee+R7
j93Gx5InOLQZzPJn7BJT9GCFmHhlln7EdP1XhCcrghRhyZsU4RXyBaPnPJ+h/xyqFuUD8EuLakn9
TZ22rHn53641SfLyDsmSSDEaagAnuKaf5B6TlcOJV+6KsRDPGyajjG/hS97nEwnR+WotxkvPdeFQ
QKzW8u/wgdSjpJvumX9F4xr0wOm/XUbzpqXNdrJ6Exkasr81/gQhMMrpGWjRL0e9gf8Kd3v7upvm
zXvZ8QhwuUocwprzMUDbGm7BsNTX/meB2eknghPkwCPOvpXMn+B/In1fhjEe6R2fJYXx2Nso0QnD
3H+P7or0bWOXEjxl6pza50b4kw0T4/IJQMUdphxnZ/3VE3Xu4ubsznaebUIEynF4+nLdm8qlEPbr
E0OAOqJYwGOtlnvkRliqe6UM7uB+DasH28/MlTtCALWA1OpumMQa+Nt0JJqpb7NKalVwKQdYpvON
RuIzE44EVhlvQk1fzRpGIozFsU3Ekax1SGQImH0umMK1h2avjVn5zP5pztS3GijkKqzKJ5dj9u8A
jO3RLBHIsCCJQkN5aRawgrI4kz6/wVUj8HJlSaSvHDWkGrugcd3b7n3fosqd6JdqyAZ70G6yKQms
b7Y0EMRJZYbLcgwmEUmACoVwlgO1Ud2G6iXX8T3ujUXQXUBGa0PIuHf4lP6QD9L1XjhBgExXpZFt
HxCcbgsZHdRli7AtAHD9z4uMwhuz9EMqCcuEaDztCamnbw6pN5sSx+1uM5GG3oLWIJrNSj5fWb8m
/XgFhmZ9/oNqgDmoz3hcw6Ij8gac+gh+tGM4MoPR6MLNuyEHvXkAAeNCMJ/oG+G7hoap3Hr+02OX
hyb+q0DSr2wQUY+lxH0v9nD8/Rc1SjgnQSNXGRoDgp53EPQwf35W2uU8PIDtKv7Tw+s/J+vYZZBf
i2flW9GCsA2ZZ9zaR0Ip+q7XAatkh0ZeScTsAn8RlP2EbCAZ6Q300t3BZR/lder9UDM3X9vAg8BS
sGXPG70gZ7qHg5tF7KWOSGH6JRjbRtuYaI1tHLuXtULlet41E/KuLkF3jI/AArNkbRX5W+BFAGJI
s4UbTkNGK50n6RQZzUgkv2zRbNBcpQ70kR47CfSbrxSGXmywLCVrb+Wiy/ZZLeKjQ2VkDvCA89V0
7kJ7Ck5hiv8rvpTBoZ73w/La0Ptv2Zpfygf4cCOUQ4Lgce3EMID8yidyjgctmH7FFrpUmXeTN3ma
bsKwR6e7/1RpGGIM+PL7FRbfj2Dv/R0RVlISJ7QrJlhchKOtuHxrHqel4Q8K3PZhcpS7my9Zi9TO
kV68tILPtPublsxG/t1P5wWPCLFucYGsaTAJS7igbJA0RaabmYzyMb0B2nTTK8MEZ3+gch8Qe91g
zOr+laAc0n+SoVt4LKF4QVLuGwjFxKb190XuvE11IsR1SmDSVLV17XhOByl8+btBe+93Umu/+X0s
F1FV/bgZ6/0kSzg46brKCdghUHJa3BY6kIaZ/E1B0Jc4jEtp90pq2PBaynIgSWooQX018pvB6GHM
M7LJg1ws7n/iB3ltgSxWLJlJu9g+ptIIUMJwywnuwdqNN071nBAC4A5CFFXfDC3fh278MD7ESpS+
wqM3q8rARo3x0nf/uQtaX1W0BRNT07MkM4dfMjXtoHn4CojZE0010xHveCABhQfjRtRrFe9QP1lA
56MTaLk7zz2VWz3iYiZm7WW6mcqMkpp0DU20vAIj9c1m6HHN0zlBf6w8nzrdDhNd6zOtzNDfG5Rk
Jl/hxzl0CLerfxQvFt5qUKXpgXqbL00SLVUIBcWZSyH5J7dizI+fJZq/0inb/dCcD4yk1MJJzVAM
i8o/Y8ltCmnhbec8TG5oYHUIVgzN834i1B3bwBmWgkeg+gHv838CuvtttRAviNpfG17yrl0H+4/c
msYH8yeOp1lF98hibEAT1mtUDPUHxB5oOm9diIdwjgEfQg6LJM3Mt8pBA0tE7i7pB4rU3uiI/EKR
Uni5LOK20rDEdm2ktMKQ8cb14taUfjGF/kZgf7+kp0gUgUCMxkNA4F3/rFOso+zUpK57hr3XSbuW
GKPWDA/I12d22HAyV6jr65JvvXXcQBGYDeefmXZ+wjR0IUtNiT8c5ji0S/TKhVeAM4NWpI//uTmT
wxo4Qcd3iLcsHfF3aFGJ5Jevpxl90I+9T/Wp6NiZmlaZHE7UdWFWWKGHXNOV0/bnEui8CStx4WOm
Z07Sl+Lk936sC55c6d7wUpcLpDFUofZg7+OyOZWQyt9RsvdGleYs9NoZDMGbv/EWSmTSuJ+QCrXB
tIxzQJelq600nkRwitQ35e4Yv8nzr6ndIQZ3sKY8aWVEwTjQijx3N9pIqvtfXcVc8d47OrldVbj8
x6nbDHLnwS40Kwu+9fl5bdiZxzCX2H+jJe9KXmF8uU54vSHYmghv6/gTE7Bpea9h3znsebLWsfvR
gvv0QXhhxZYzOLG/K7v4b7f7P25CMDHs/vD+ysYUD8mRhONFv7oXRNwLziLt7fO6KjhnHhQ/rk9v
ig9mjZC9PaPHM7xY/iYsEU68qbaYUTdiBRUsS5lFz9dD9SjulrJJrcFC6v63i3d3CtvQ25ibNhyj
R3hCr05YiNgwrASOS2DzQOjYht+h7ZvVYCj4HSy7ghKLEwzXviSGqAXUFd9ba5g/Bk2K4X+oqCL3
URcWlD787eqBTfLP9uWi7p3Kv4QsN6SSBsXh1V+fdNDdD6hrB4g13YGzIMC4mZbidT7LWHwfH2Km
Dvj+mol3MhboOl6Q95KftPPlzo6XbPGsPJYh/TQ2Yr70jR8qCpGVcykqNm+8SBiU6OoH7cpw2t6B
TVI+W8kQjUj7TkgzASZuKeo6A2K3nUBBw6ykMIcF0E6F0qWqfO7HZqjR4kRxhO01FFBVOJpN6FHB
Pibd2f6yaLjECiaxpQET5YC1a4kQjvH7DfEn+YsViT9lHi6WaVjyc7x924m5K44rcaitp9FUI7+N
uS/T2j8iyMvSc3LgtznMWEJEdCHdfkJHs0eqEFyY/yKSLjSahvJ/MJ2SLBmrYMX9Xxsn7akg+tyS
nI3JtOPZGSIAxZE6igrDkUGJ4eifM9CWn12wQwn+Oo1CGj34s9TwBe4H6vy4FYfuAJ/4TIi93ekU
cJXBzLassKW7rUqmfhRshsfoqBPhVGS2aeUiUgup5jyTXzs93S+F5rarUfEm5fDKmBbs3ByDe/d2
YWpSYiGOsGbTFf5EGbzKlp8el+L0g7kjByslerC59tl/e3xRAUM+aHae/Xzd7phVthTLEvY3+3EX
BXTVidUpQ09S7kRDLR9KjWFm5RVWe78YF/DjxXVE9wUSQGMIpJYc9E5K27fSvT96TIsEq898yRf/
CvNZapH2uE/vulgPLiTSODr00w7ocO40zVeXQZna3MJuf7XwQrRGMFU1FNqgWofHrrVeSCRfqNcy
FJVn8YNhDMFDuilsipRoqp/3zM8ZCIpTA7JtyYfvxK+WOXGKgc88jX57VneGu5RXVaG/Pc89P/Er
tl0s3csSM0EvHc8QMWYY5W0UX9MWLfF4E6XD1LC7k7VxwVEL2Utbj/9EeRc+RCg47xjv5GM7CCd9
QEMFlZpUVIe8lD5YxlMCssZ+7W+R2SpJs6gmmnM4lCGPrAHutxEBRSpbCFk3z/7uoZ3JgVv09agt
69aK9j9gbR9E4xSzrUCEsdJkPFztcWH1ZvVXxj3bPZzx1zSRMuuhuOMtLgusLwU8Yt2p7qjK9Hjx
dCr+B7rDTtOiM4w1ZBOJySTd9hwnjxY3QzlDaJvpUisPvwux1w/SqCt0lkhEo6Yu5fE/xh4YoDJ5
OYltlKXeshIe+/F4JaDIHvPdRcADjBenTB7gz9pwOesgV3NjHc5QaS+BXigiteAlJ744ZLx4a9wp
OGiDmoeQ878y7a0hnxdV1Ap2GIEbr2DEXfnTn32Bd3xZggCeabMN3ep9EdaS11uIkkX/RZmoND6R
ssdT/sZoMvxoErz+oAKTNtz1g4yAAE1EW4lyeoqfSUW3nUOUZwm9Ms86DHffwVcdPvUPx29fgoUX
pgOO0PQTenOdF+104G9Y2rsa92tVZcGKm1cpUgCQcDGmP7sW0Nl/1IwvlSmJtQLKuxeshd1rjmjX
9TlqOljmbYTV7GZdSYNdG3k/C+k5GpBf3v43pnaD047lhNicwFv0dOzSj/EglM4+cIppx85MFEeH
mTWpo824Kz8n8AwchB1SlEGTWvSB6b7Te8LKLbm+DqTP+86ALx+84l9YieO2P5BGzP+ZUU1uuY3n
EfpsuPJTXdLk0Kbs/8zUO64YaGsPcEAwPNLV4i2s6gkpTC53VvRtlNDIirI75K5K9omyFNlGTc6e
lR8bItZ8Cx3plKssxe8CeKrfP4cLCf0PEnnEtzRTJcHR4oM9FblobmWr4u52pFaQGjDgWOhhM8Jj
XliPfg7ScdyHlJlVXDO0dNF7VOMqrsjEfLnsdYdMPuFG0i28UdGFpCncVewmpyYpUff8cMATpyDF
gdhrsUpo8zqtoo4GLAmfEvzz6LkTKcgakH7ucziyOtOv8T3NnfXMOlvTVnTrrKYMQYt/XVFmOXFo
cJp1Cmp9sCmjbIFhyCAUet+zupL9fnsqCc52nykt0Elaq9Jvl/t20Pi+6T0rBzwkW95RpDJHX5ZL
nxryCY87O2nMvzrnuCDpiMOCTnDskgVis0oaPNgJvlSZbiFFe00/0GHfqqR9Xk4bVvVi+bTTTwpn
OJbnShd/jyftSiBLt6hkhz0n8BZeQrX5SfcHlEu14efqripn/D5BqMOEUDeY2DGZ5rYNJGuS3X3A
McBAMxJBQjgByWXTEBw0Fof+co6yBUJsjNt0DfzixBwzgm4zsstish4vmfT85IHltC0F4lUm2ZWq
tYxBjRLhOEZxPRyTiqMKKI004rrjF3LgJhf66bfDsyrVwhcDT8TcDZPw10m4z1GajaB88Jx6luhK
bjhr8bm+X/UH4gBG3Mx9tPtW+bh8kAC/Jrt0wjd4JSKSqpGoEbNhZOryfgdIQ2NvNV1MIjN1NVwd
gRdkT6usjopCbMPNu7S48T/5rG+BePv4xklxHSiwDaCWnYeVWi87tU2zaR7u7uOsANZQA7KL/A8E
3Xg0QITf3RKldiO7UihAFiy00v28dchXfWnlIQmKYAxNRRdcG0z4V/qmlnapffYQpq6/Mt/brClk
cMvdNgTyXzD1ED3TfXVc3S58wqou5YauZ5VnGdJJjYybkF5SlauMpe9mS3Ra7gtmJGsHHq7mVMxb
7/F5pwr28uIGf/kBtlnkQPCFXRe8myyN/hD6dPCO5JXyoeSOtOzhdMjrCkTdh0pLBvP+jmZC7spM
BIt0NHq1aZW11yDz3AcdQNL+Hvpu0F6VYCcOdzeMkzD07NsHG0K3Vpo3fQBUXkQymwqRJnysleE9
WfhBPjK0auw3mWZNOgcv8CHu0hpLaONXkISPOl6aMxsMBIb7mQpZ7VvgLbQ1PsWeCkf3gnWd5AMr
8CHGyYcynaxC6T4ybGD2eEF8um9mbONb7crI+2GewJSif/sPDQxCwoJF503jlf8Waupx6TT59uvv
AohOYTv8JZqVWp/BeM9B9/hCENteH00xBjqoU0bRnxTe/MIjen421GZ+ZnZKZXciZpJE621/0yml
ia3I28fFJ1BS0UUG+5Nq+oTC2FOD/EO0/GdPDNh7Dwvx48HP+Sg2Jypxt/sNJ8Z90OJT81gMhgRs
0L0kI2hsrsmD+Pxb/3l/LbhQCGZi+idYix87o5CoM0HGmejcfRgMOzihSavDmahs/7tWkcLD+JE0
lIaJ1dRrhCghdCP6TBECtpW6r/lC97n0GshUi0IO8SfKHCxpix8kqll3fAcYbMhU+XqvS8QvuKZs
s9lwIjmM7tWF0Vd7TMr8ioP20kwj9Ose6SbsStv8i2lytH7WpbU6w2wCr1ZnO4zFFO+mTpcYJY9y
ReuYaB4iUwrnURA744Vusg/wyOgO78TLuvvTsoZssY71L04C1dHSSm3oFqq51rY0wUPeMENB66HD
C1iNAZ+sVwsuoOf/N6uvyABwKFk54kkTbiDRDCAlhea9i/U38jBAs67WLJHHqpwVWs0PosIjGlb3
gd9fIrc14q7XX82ccbtSitaMf/VgBP/RhGsNv5QLbK8CtDFdC7ilgC+Y5Sz76+EW8SGynXAut9gU
6VfXaZUFrKTn9zyoYbZKMYofM55vTDyQrUnu9lkVOUM/GpyKL/jTCaIkEh+akH0X+H+oFGsBV/EY
HdzZtbrybyrOCE+Ki3vaw3gABQdShsFhB4blg4MQSsES4AVQxr3RWU1fmV732AIVy3BOHJmzXqCs
Ba+xXk8oJkiPAExaRsxeTHJFDMVuPgPsyncyFsKuGxZHFDSQEHoZwb5B26hK9L4DhBcsjSe5SPkr
yQLTSzH52reOUqSMmkQeVJ9ld9XUQR0Ds+4+dbEto/OGgJOp9wEQR1njU/Q9kNSNmE2tLt48M/WJ
E6D4wXDJ4R/mJic93kS+spf/W86qmW4u0AmoPHfejeGiGsEg1XHmWDQVpwg2jzR1+o2SX/Xu3vNf
sOZzxXJCiESEsk9Jd1DEcd+2yFwfzJAoAtCdaMfmVy0KiJVA4DJuT7zp/hrIePtvPwXL9HTCoR3S
6NNQeCPAcQlFVFsE2m623IiDbLudaIsZuwQuaOXY1ls4e6C21Md2m2RoeDXH3fNKKrTg9pxKHEkS
dMSAMpcwm/x9zt8P/TYsKXTAW0yluEbXPxOUZTaqk7odnkdtIM6kzr/4BLFs23BEpIpbMzVNZjsk
8mJdZoOt1AL+lWsuwMh0aCumZ10i01usVpQH4XMeOlHNX7reTNELHn5/AjfsVVpuG6WMH0OnRY9P
tdtXwX2Sx+WY41uK2C1Hs51eU6HEBqLaWfYpSv5RWjT3R2BhijxnRGDzu9LY9POjgU8Qdw3q7ctg
IWYOvLL0mwAhebg0oRTqcr4UAQKqI3+Ccnb/UM1sjK5u8B2FQs/PwbxzaftLuZjOQGF5n+0MP+wF
dihLNggMiT3IWvJdQiGFMfcNnIUsfxToXlEvpi7EjW1g8IuAJ2rA9NSyFUY8icFtcAFxkB2y0P1P
OZZsAXk87QYDSf8KzYW9JFpk5b8luPgHpwXa840o7Zq9Nh6cSE9Zn42ZprgnB2idcsCCEptn1HeK
pcY9YQsIFsGeQ6gvQn4h0/N9hVhEtlhPdSiITDXO3FxRig9fnztR7K8hX/C9fQTOZgM/rPEHnH/o
7Jedu1GJJSSGqKPbAdXWX3s79/mDsbZfg0fJiQR5mes5BfkMS6kt8raLnbaaQ7xGm9uAoJN9zr1h
0NyD2no79juyE08QPFrxVdO7BOLLMrtVJ/Zfw0fu9FIjX3zlA66OahDiXEuzKEwj0vrMucz4Mvfi
WSOyruB9/hX6peXGTIsLHXRVuolMdMGkCh9Ce80AFgzz9AmfqfZruQb1QiXNQfDnB17enmuOqNAr
c9Zxel6L3tqqPvWb3gcp8MCsNKr6VHMJQm8rCOMgZmbLNysnfCAn5y8q+lfAYoKtRtCqklsZ7NM8
7mteufohGAWQ7ugVXu4qr6EbSNTaBjwFTmkC3+6+/qnf53bBQ8LpQpccMJd+wICOFtChT3N1e9EQ
v6aiYbudUwOAVDVQIkabjwN5UDCC741iRhhAePAG4nETiommOk3CJwAQhBcebtHD9makxeS5YcRs
SmOuH4s5QT+WpLB43STEF/u8SZRKMpy4EoIjLyS2rydf4nkWCQf9EXoFwk+ZtNlxLNZQjDEa26yu
IG8m0J2itaPfogSyTFwky+TasehO1k6Pi/3WoyWJ+IUwlJ5G2XLfvXDNLiV5S9EeIBeBhr0B4Xtn
a11inO9b9MlyNiwpMhYvK58hFiRYfrsAUFp3TJ7MKdolz0Nply10Ss/JOfDnQyKqxshiHbnk4O24
bRqjqXYlgaLMlBhOMxJ8bJWVCiBX15dV/7iKViZItSJh/ZnxtWCzXBwmwD7c7oAKAjf+Y3CSSJeh
0XIXqYht0PbDs8wqTjAgbqRdbzUJlbZ5rM0D388W9u8aNL1PBz/EcE2/8J7amcd1wF0fJo078/Rh
o1thN0kg7P5wS6bZ1s9KckeI42N/KwEfag1KpurF7KnK2CJ9qgQ3xewR7/iuGljYgSBvSDY0OPLU
s2z40DL6k/gluKS3IgfzkyCL3VguP3XHZ0LuqJ8XUaE/nOuhDFrm+r4byc2O/kSrgbHU4FK6EPPs
Zc+/EdCc2TuS6VOyUHjdnRc/ib/P9aQ0NkVFKvYxK12uX7Ozgc6PCADD8TfQTrLVqA8XcAFV2je3
sDW6lY5kmoXoC+OfiDp2ryS8TI39D0J2MMUOPCXY6mQmr9zxIcKC62U+MwORXE9/WUM5R7+oXzm2
aTyHFzXzGqhlOALnWIla2pkDIBC0CShhIM0EeTSqBk0Q6qzi8gjTl/PA0I+6izQPGnji8dGdq7AN
pXG+XB2+OF00EccRyXr8FgjUBgGW1cqdmD1DWktUA2NG+ccf7oWSjf1LVOnzwqPrez9Yr1tCVvl6
qt7tJ/sT9vMXQniE5iBo1Ajo2yrpLNxE+z2eqHFXzkSrOWCoXs4bCF6b0d1l3hgvqlIqgoiZsde7
OUzbrhtbCsj8ITM6ha/tcc0bmTW/FAomcYBpEwMJZabET0eTwjiuiHo+C0HL/zwkunCh5U+g9IFo
Rr+Zd9MSVQdNqJPyG3W0PcDYDYw2FM6Ket0RyQa4y0ARSU8TwsQubxVyl9JEHyso1lEdE1Csb4q8
H/Ma/ZSEQ52i/KBe5vYI+pe2yGBsklS486CmBnG4M9BSRJ3AmH2RQUxBRm0bfF1YoH4ycr3xny6U
gV+2CHXEkK+sPnzTjC3tHiEyiHeh4kQ2v/32vdLv1csUSjADBsUagTLoW1yKVyJjeURCVvu3VyXj
j2xZf20EHmdCaE3FzNUS5pV105FdpK+Tkg6RN0r2seApL9yUltVJ4qQZ8hX0rHjjEX9siTWR94wA
brUkK+JlsGDnyEnnAmV8VaK+VOiI+2Ck3K1bYC26iVBiZDwvo6/sY36Nt5/UgpDJauGzHODdJToW
u4T+LK/PRH83g1JZjBvc8Y4nW4WY93vWU+In6g4ny0Xk+hQQG344+K6+wUTuNO8amOPxAg3YcwlR
ViG2/iaNCpI9IlsnMB8IiP8dhtfvVb/EJwQnbzuN2x/P0uMuTQoNs+Jsrkem/BiDcTaMe8i1kJFd
4udb76AALg1IGMrGUnOxjwvkskM4Eu66S3sg91wemtbIr/7/ZsZMq3aT3qw31q9TH6mTjTMVDSZT
Uno6keYiT9qdBbbbbIAcKa7kKgq00UuGlIbRJ3F61wwL1AYsSs0++stnJiLj1XGKubHtwp3DurCr
nm+i7xLKzwkvvl50BsSdCp908j3c65hT658zSy/XHRFVTouAgGhdeH5is+MxYnqgisBwcla4eSJ0
4lxl9iPPWinaGmMJdTshI2MUNQ4HCR6CDtmPRVjc5jfq9i05euSS4gZeaALB26hihA34Vo+d+T0S
hmY7Fvo4VRjemvEQf0BB8G9oqwMJCgatACr0sv62hPEvC99+GUWsVA5zeDzUrKbz7yanwtBGI4on
vC8HS3tU+IyKbmyoRPhX0WXp4EUUTLY5HfnR+385MjhLXx2dRBbpWoT7CDJRIqdJ+i9U4KFdYBL0
NTY9QuuzalhJFi4H4SaSpfDqFxwrHfoMXdLYejNlZWWV9Fxcdiz6347BMAgMmSo+pzX4EnmruLWK
SRBzmTRMIS+E7s4inmlxoagCda7hwdyzql8DcszpTFI9NjXNyChaRtRYWFOfzE1d1zZIfhrLWqzp
9CTsvlAxWQfhplIDFioXJIsQ4Ys+FWRIRLiDybjf+zjfYoSpORxNWJzr3O7KXnUST6/utK1mUnQV
rHDbx4ztWkfgiQWo1u0MlQ/aNl5BFre1xSh57tlJzVe1RAU1iOzdrxmUNPgjAu2hra2I/OKvWUMr
RI4rjblTdAPlKVtdsQ0gGTRG90SRtUoT6C8JKLKdKF87fFHhEPcAt2QMv+1BuDzPxkmXX1F1OaIy
I0lwiNeEQuQH88WsTWF98ilRLYANqEnyQfYYbFdc98YyyvjL0C7XJQXr2Lh+h5kxP/L0ECjsJquS
JKVSs5r8CGfrJZZO2Z0zux2AQFsBtNFndGKFcV+Djb0pe2CFhsg0+5BtLE2gcAudXdVt5iyavBfi
ACIDvPSGbZ/M0U3t9KoRUy5+EnWTeEUNF/adyqXcc9M4PrDwi1BQ6qS0F5Qg+TsbHEuJ91FksVTz
yWjcgpVbyY1g4bKAMTwNai+MMRBGzqaafC5uVbhkjLcMQ9ndYg3pka87oevjtO3jLkiJFQaFJsOv
bJQxihoXb9T85WQq4uixwdcsXvi6SMZhExvBmNdpAOpRWozv7OujgUSiTBgMZs/MFvmKGdOAwKIO
N8CbFlEpuANM2YReKcd71+p2aHmXi1ugZDrV5eI2GsT1hqO19JRym3LTrdnkXrBPpxVIFGdGtxQw
XXlZheN6lseoAgzVMj/Yj4XYzv6+o5g9NMgiWKI/6dH3bx8eFhJ44cITm1vpAlb33WuUbiZD3dBw
8dShFpwwFDDNUFQKPruDJ6dfiEZwnv2f9UmmX0Ogb13QpeQVpAfBuBnxf9Zz1lSeJTzvtQJwYh08
tbNX1UVnxJgpwX/mjRRzCDJflVO4fi6YT7SHCfFTbgot861MfotZcjluW/H6TqeNE/hgxCVIT3RU
nDldpLiQvwKconIDCdLuBziDb/C5330iO0SRzyn3ldmGUUq/gVwWi0wpRMa5oxPbIadgrEs1jUpD
NdWnHtD7uWk7aQH77rgPfuivTaLkWVjtGwBMbx1MQwXgROjwb9ovQhuampGm1Bu+8Gmz/DE7kJO7
Zqv+eAUnMHxe1r9HDUX55x0ErQ0wiya5/49JlZJnofOssq5z4A/1XwXoHj6z5Lx+KGvJiu2nZycH
Cs6rgZDEFeMyqjIQFjW0gDUFSfON5hYwGioyddyPQW8eN+VPCL9axKNQC8bxaJpwTlx69KEVnnTW
sPYvRuxLvNz1nGoJeWf0gAN5t7MGHo1aQ/P/exfFkzuHX4yHwmOwFSUG+u2MoT2iZKIzqx5pmUq3
FjhfSDeo4D+HsTm+gvQ7UAuCtYm+6ydJD+4bxV/z4R57Hq0n8w7wJJszfCwXLTnpFq507E8qVoRY
URXmvBASaKFVDJeQbKTQDk5LZ0Ivmg6LmeTJ7XLWh+E5BLlItL/mDRCjDtQ9oga3dlwEAbtYUXLi
KQ104G/i5vId8yO5sKqYh5NF2Sg6PDjimBk8QfplQzxrd9px+8kqPSu85s+8pSk5/lVPige36Gqq
byBnRYGl4cVBrbHRT8gy3b5HQdImhQdEV/KkPIcHJhzHW/OVlxQta/NPNa1L2Dh9xEK44ZsuYGEd
A76INM/65hcvFbDnb6T2M765Nvi9TwkyrZQyfq/0EpAfKJ1FDXDxbHVVHUjiUIDojAvDh5HkisdQ
ReYFKL9PaaVYET69JamcaYYHVAWDeaVxOsuW/VrX4qshThUWsn6DYzOp70GCn67vsuk2uhK82Iyk
D1hNfGZ1G9vjS00JjihoXoKWMVdLTjDogU5HubQumAex8RkBMV1Z6PMGmp7Nw2RgIs9+12sGGV3A
dGGMtMoNcGfgiaasew69kw/Z4Q07oQEkH8/oW+dS5H7zNcFSMYM8lTYk8sNGsRkcz/0KZpIaDYij
ltrw3Ejc62+TxMR7m/JoyKXXXzpCZYkv2ANxtA/9Gk1L+C+5lcGvz0wHEgTWSMsztU7Rf59MRhmM
+U+6JcnDOF3KwzEFLWZk1z93+Aar01/aj1p/ta0sVzNzpIbaxLm3mP2jCs29lUGgg/Vtu2AdzuCf
DdR7+jIGuOOyFZxXpZoYvyN1XpGeUrD6HRX6d1JiJAzzctlXwo/FwZsZN+9IEuywy1pUDSIVmc8V
KOi/B7TtXOsi+poodHqueHo261qpQnrTQwA2tRL4TJqOn1CI3RGJohfq2TTf18fwzHOisCWBvnlB
WnElV6B+H3TgY0KnSXH8QxijzzeZuOACOITJNx/8VrLSO+AcCTUKFxuinqVRUYOxRiSf5CnuRt+5
MxdZDbmFRRCZDLeVqFgkDeoIGxm6cMisLzpojczgZ3q1AjX+h2cZohb2lT68CjtgYR1izy6kjJ1P
4BR3TZvATXZyfRUOc0JCU33eQUQerkwjX7yAQ657XESM+zUa4tHfmHz93fC1Bo2XX+Hzy8Nl3D4I
LyWjDzvoGrl/2mhh4SAKiLu+whgQELZQ6XWtlMPsPRmk5znvVG7BXK9JtO+tULRU3VmRdIwisEpM
ICSn1rezYzbXTds8nB+eZ61goIKjCZcstxwAz7ag4XWMnIDE2AVnYrz4s9VXSjvhpgRowRF64Mv2
uSJnSuO0Aj8eRz4LJZoUx3I/IaEpSC7k8X2SDtWgUIIA1cUTOmtISGQ0v+FDPXuftH/Pz4S7WS5I
aw2JbLLvYJ/KPLyKIVxxXKOPZiN4JiY99NTCZHoIQPyq7w7PTAVNyYHC1MxQpZL6H6j1cuo5Ebgo
Nj0Va6+UkTntHO2oA3pNKOEGnYQyiI0puQCQF8NG2gyz6yepqq6E7+v2nXO19J63oyJN+p/jEv9F
hSrHV4A4/SuV44g2kFLF4UvBVaPEgOGrjsGuERm4nXRcCuKOvIr+0tfTcfUimT8Hxu77TNiCv5AF
gyDKfhf3rIefsuM2ZpfNTSYO1h9uu9G+IMcHHZAIo4zZp90oYLv9Nh+UQObi5JeLduRzjbIPLHuj
ifiRKd65xaFBGc7fuVGuMTi6dWvSEMD9BDecJ4zsrzx3rkJn6g2E9gRlKdPOdnjyDjKTY6Q+gyzo
AxnonZsNVJbvl33w/BRUFWL7Az/P3BAU1eHlUKTh2Bq6i0iyRIvGazg9J6HirPS7/b86K8ux6OIe
6JMcCiYHo2mp04zSlrlxc5WzjS9O59r/hZqCG7Wlw/4TAQcsy/wd7kwjRM8akI7abe1OSYPeYE7i
aaU6VdSv04gfIol9rptgCNmDOY6WbZF+J48OrVNwuGkkKXGZw1F/Kxm8d3rTQAPajCRIwzZVEHoK
SFZ/MsrYnOMDTbs0ATTjD33Fwh2dxN2eeuhZC+Lc0DhqXQZ80gnclrG+KhAtuFlMIKUPRPALlrjX
s1BN8QA109yoHtG4xKrAKSp31jk7xZDz/MUAucGojRAomunjtfO6EKF5vB6mB1L9VcAzjenr53jN
kXSJZHjLj1z7FqP53R5Fawx2dW+xk+kJRx4pNXbj6VcQArYVJ41qK0mnfSY1yEZYtZD+xlnfDAaz
RgPEHGXh1blZ2AEDzUYKJ1Cmx7oAZllRcqPvQaZyCfn6yUB0y7YpvlBYEAQHfRnfswqPDhkArLH2
m8ZNYA9zRKAWS6K1pWdo1lArHtpiI5DNriAKOhRRjVKKAEeD+fr3KTyoFqZwvuz8CiPzDb9gM2AC
aSZAq8F5MEIz2b7GbKiLB8psblJNEYTTboNbScl84c1pfV+I1Vd60Asv3tUwAbrIRFfJWLA8ULtq
YqdKNrHCFhjP9XxCZGVBP9PtrnZuzjvdaFBeuen/O4QU5d17ffX+JanScNrt9teJ/YuQY8CkuOgA
XxOsyfGK7ElFpp+YY2UTGrx+QbeWNs24Z0uRbLDTkvwj89CAlPbWcBmOnkhRc1uGWJRkoBvtOQAd
Kmxz0kxa6sXdev66mN6qRf4eWc0jdo14vVZ2xsDxCs3ATimKIlV1at38DqdGVJykGxzWBKR/ZpzC
CwyCXQi1SpHmc43O5BKBLrBvlHbQZ9EvmgaVGa1wYMI9d5Avu+iiDgXQfNpH7JmEm8taIqWbKvb3
TjmSv/GWQNCo/KYv5Gudh6J5aEuurI8Tz/olZU6RznYKbOGJjGAZD7tcTGRcW/oVFcN+LVZUEHNF
MTj1+cTTdByV7Kzuo0sbM5ka12DSvj9GOZG5WbmEAXyXmMognZDSXXy6g3aacVqs+VL3/RgVpN0p
u1cG8HXKoEtBYTPhBH842Sv/vxbLUcuUweSTpAIaS5QXrDRR/1GgWiqMVx7cXKOSanSmTSryLbWZ
JB2eVAszfhzrK5DWgxpgbwUt8XHDCh/hWXvz/zjrez+NEXuYFbBynpHkASdXzBWqHw8ecbIItIyf
44p9UZ5uebzCL2Y2Sunx3WEMOZ+x81M/MZGyDyCewMzcBe90Y/ZvFxvgmW3gqDeVF7+fVr13f5pm
7DlVQV+BgRl/6DRmCzUJ4Ukwm0Gcbh3aJw48mp6CCaluuMcIYXaof5Ik55KiGjqEfY6oSL/blWxk
dSBbQBEsM1fzxiljLKrEMIMvfB83GZXcW8sbHmu2h45JLA8t9vDuGvQU1oTN5VKZAiXuPJeSKzVN
GnN88N5kCdUXwBIvTHSpjrVZo2EItCi1BVryIMPbiFJhrq9X2golhYojVSiOf/tfo/A0f3MNzbbu
QwSKmlHNwVd3z+/pz94u5lOiXYGqJteymPchmNZa20WDWtHLdNDAyRv4by9waiX7vu6UaUL4XEBc
oXI+uRICUHO+yDghBR5JNX3idWf5Y0IFg8lQCTbgbvBLC2Y/BaHaCLlegxi3bcG2pY8xvMA6TV7k
rr2vw+OtggO3FANzvW95QMVDudyu45LYRu6+CKDTJZsEiXZn+22N1IMD17kMsowpDLbVW55gobya
4irqnQsU5Z/IUXNTOdi/TLd1xTt7YN906sXbf1mjRov6rrPJRvS9oJhMqKHBfdwnxqqPy0fnkJya
aC21X2TY0zLsuSWJFLQZJWYnSFvJXBDRrySp7Q7GqPHHNF6QOdzrQiVC6hxZcPwWFOLmMaNXJWqe
sLWmInbiV7Ncr0eVX7a9BzK0YEvvxRD4JRpkcEdrD9MMJxJObWHVLZEriUOvTY9F/wreEzT2IfrS
4+VccoGL+Rx2Lc55lrqIva/LyxmfpXDvyUJqhEkOZRSKzVaqPI+LD5C/04+XbIfa9CAYv/PYvn0n
SYonBGNzldI7Ym7J3ikAEgDqtd78r6xDB2KrLD98EdJJ1l3DrDtYWhVO6wjP8E3zAM0Mh3Ip2pcW
Ur3fkuFLLYmV6gNZr81jguIpKPlQIvuvel+Zx0g7bhmmRS1x+bRmFmlWYhD8iVkkOniwSPA09vJf
WXWfYCGlCLpsq2dlQCgjMpqfOdxLVhOROAs1vR338idlUena9sOgjwJt7ySN7/ZnFAfsvRTdnnaa
k+4xwzG11x2/2F/q6gTrLTMzzQ+jsUVHpMFTWN76PWVoOLrsL9tWlKtBjavzyiKzPOVWR3Ppx+qy
nYEHypYYV2pjMmEkFj2TY5v7/4blx832+msNQcrQzhzZZ4ZfzSz1bRuCrcLcSgApzgf3loueopDh
c+XpORiQcIwZYwogqNxosi9F158mmtw64Zg+qVSrJgwTWBodXUhfRIwBLk205YwbX/15AzFRg+aR
2Ae39uXHWKBCgjJLHkO7B2VT/EhPM3IylVb5NUyuaeGW07RwX4gFjgZKljeARpKF6htF5QCu7z/i
41rWdd0ga0CiRycjTMGwP7KaPNU/amlwGahR/C8C/4/AAJ1JtHm5h6QiuJLPNXocrMmy1lYgNpQo
iTh+fjJ/24orqFvu2zgFc9LIATCzyAlDTwjW2kXqvkrnkEgZC6KOQ/ewk+nSPsB6GwvfHrduUm0v
AFDrhmaz8AplTWBqQNnVrgnoX+k7yVTyD+2lSRJTrjsoZgTdQSogrXzDad6blZanb74g2rTVeSEp
5bR7OxB+TG8k4dEFhFL376/bc2Y8afnM2qBXDrV8psaC24oJSSHg2skU/g2G0OrhV+C1NY82Sbth
oOO5+zb+15sHKEDyo7f3MK9Z27/f1tsqhGHHVLaH2HWHYIk+qzTarNOtlU0wwFaNc5HwML9I7jtd
oTnkMemgBOX0CkytPJChopVwoiUxc3dbgx6tSN2mhq6bhNAp/UdxC6w4VoRjDAF3LH+Gtgb2dX6h
nnmNF6maWtAzJwbSan/MqFxAkFliKvpwHTk1d6aSyVW00WlkmxI6tQUVfGVOuEOAgXNUA05XHAx+
hkiQZA6BQ+RsRo02xTT9y8f/gsRf1/Y/jmgAUyhWKW4G1/X4JtE2TfwQ4/eISbqhughpYi9kIKRR
Hvo5ZWefcy40OlJo0QMzz28KmowtLvuQoTzq1rHjM/UtWc2yI1EJ63m+aXj07IwCeFUH/nS9bx4l
Y0QSx9k+jeVr5OyCrS2+ZMtWmUaup+M1yoRM82PnEJlTQqi3sgiaQJ4cPPlH91AgULk9QP/6YWiT
AXb7T8PIfYnNLOv4LpJ/HMyvkEMh6Owj83izVYtgGa+iDm3i4VYpXemVBJziD1nMjSRWU9CRqFN0
jCUKuhkmXJ+uN8ZvJKRqxLToCFn6kSQKlhpup0uFXDlIA34tCnI22pKcnK/rmBwwPVUpRkNGyXiB
03YL69QYItT68MAQi4bWhBErbudPxcPpHm3BsUWuqQInVI7v6Rx5htRoJFFFBBfM/FvVVo2ncp8j
OWNZ6ednriCVXgdGCSMqkmJSPIIrRiJy7LpS+x6dWqSegxV39WBUmYzdt1cs8bwRAY6MqI/itMH6
SzCyHYAB+Pgq1ZE4m4cFF/UQr7QV6VtlSqnXxBTWNATbVpg0TWfAJ1Hs0azcz4lZZY7WqGqn6OcE
sUACpFaXliNmBLd1dyDr9xSdpEkzctNuZ/vEFNXKKTUoP2/+CjuQhGSe0IKNbZxXyOySRV8bhoyG
0hAEv13V0F5CLw0ru/4YNM5IjLAx2gzSq6DJugx3bSa7R7Ukkl2g0xb7KDlxlGEQyLfm5uy/49cH
JkqLbWZMwu+w51wOJWTL4Q1S+kaLTDlLCh3VurItHht/rxENeG5yI+iDoHDDm971nUFtSZ0j8awn
gzU/XHP0gMXwt/3IvkjFDyqXvELS1yz9KBpoqe8A7E30bMdA/ZQC6sLbSxkXn1aCcLzIdmFIUsc2
2rEOYn31h3D/OYuQKQmyt0cH+n6qMauUlxYm9n65duOcsU3hKeXFciB9bboa3VGUOef+KH1kNJ38
uQS3K+BUL4J3bggA+b0e7/2tlAlBkOk1enFB5RhNCj7sEJ6B+lc/SGGMQmCbWC0z4zMjwMgxIPax
lQojNEeIErDaa2wTnUyqMKTZ+3L4wmDrfcnXIXPYq5GGCVzoGh9N7l1RwuSvL7EMauruqVZ32emE
vBMQgKm0Iu7f+rNA5EgPCat8+zVSBW2JdgyjHiZFyI8BOKSEE0cWVZeETwHL/cxBC+8XX9u7HqTb
f+oiGDE9yx+NNhKquSqksNBgp5AF/QLjJ9/xHmKwbsF7y/Dcqo5ovncJZYJ6UYT+Hv4/2gFYt+fp
p/XLyBI4x0O8CAGken4PBtqwnqVEb5rgMV4hox8WNSMLgr6MH4TDABWC9S9e0U+KUiUXu4lhY+fF
EJ1B+p3gm+6EeRtmuk6ywdd7PuX6RmW4h75OFteCHogpGEJYRcWLx6oUOVA/Ld7pY4TMGFXix4Gd
G1USGprhw5R5T67Liqw7e9GbhnJI1kSOG3C+9Tl8V404E+0fj3OpNs7UQtpJ3amcE9HD41oXidYF
UNRYbm1kfFb4OIXKPDKoY0Z08qlSZIJ+81koBZTIBMIsiGTRup7UmBDjQcCYI/bl1TkY5o2kFls/
WTYmEXiQMyggMMapyQaO0c6LwPYMPWKNcJRCHXXXlDQ8aioiSvYqQgSpg1Lzmn3T0ade3XtaURT/
iatH5Wgiilx5DJZwg9H6AFflI/OWUIPR0c4XdklSw4UrTKy4E4cV/4Jlfb18CsEc2Buj/1vpezCU
KGcSdi52XU7Z+aU/ic9v/opz8rxQVwIlthGAAhka0NUc6K7jNF3lo6w9mcaLNLsLsULnlNpAApMA
GGuYNMZvZNw4lznn2zK0Fvcbc1MIiQcQttCd+ACPjyV7vKnI7lB43L+IttTaVKv1EqWfzhp5clQS
gRFker+tDYZ2HYdrOj87z9yTaEblaEqcTOoDHmz0iZzmlIC7KUqlGSJoxcVjHAdQe5XjxcE8u8UI
V0C7viH/pwAGKHSBYOh5FexwlEeKJiBmnPEvL/NqZyorEG5y9mMiOTe0eV5rSE+7Gv3DZoHXViMd
LhTg+5DYeoeYvbY0ZhSsygno4+65FoXBNfKOKY5/XHFEywdDOG3qrt53bA7Hl/8/h2x1QXeTSYsf
NrHGfQAV1lrhv7tod1I0ehUs3bZDLEHCl2Vcpp6CcDT/AV7R28zZ55W61bTIasggwPCRwvnE4G//
riMiEpGT4yfuYchxVVAKWCABSoOoLLIwj7eqdavM7znSW8W0JM1wl40fBAI4lntWioNnLICfjlFi
usNp7waDDBkUNl+prCfYO3av3wgu1MVeZKLVokoIQlBqKL1pjhwmcDw1BEi8FRXb/Yc6JgJ2VNnQ
ozdRWZZ7rCcVIO0BDu4RGiIkNzduTPq/K+NJOp9+91aJ7ptr+zNvO7/M/8uZk/ZGQ6ruTvFWeXOr
Xh2SdCrTUdd4XlOx7hulKtMkbiji6xKbZuKURMORs60zGjYTw2Txilx/seR9Z5RYMNpbnuEQol9T
i5uN63k8Zn3ZdV+nfzdh8pcYYLzc0msG5ZFunUBZIkh6VYYtQ/QDDXWWcO6mLWviK3iTLm71wZ/7
//Of3U84N0EyA+GFTiDOnfG5lI3UuWa4rrZN+WWmRiv8QuxLS64c0cs7nknauOR2qnA1LW3lvBQ1
yan3mYjx2I9XckB6iTucS4gNDkneWNO6kn9zvafe+P4dF+LS6ufPsCTrMOTwPYuqzsrXVSSjPAB1
+1E3YyVt2X0of21TUCC/u1N11zEcW7Xi9CUll0bfjffqkWphJNOh04penZrDP+omeqE+ZpYkSYhU
1hJBiyRr9xMQsRFUTO6uoEjUmeQgg+KrZVQr7kTcUkE6DicogKR6MoPOfZtE2TXmNoXUkCGgqA3A
s5ODbbDhPYVM4Q0lqsCvVpLIiI4Nkt/tzgTq5NnnuIqWXQCMPWq8TLsj1pYd5x3HTHD18ePamgqm
aHRJdUaxlSuZyluM7xDlyA5vznNrX+in3qZ8litX/soKzTAr1FLyAR611qVlTNG4ld1yo5n+NnIp
zRXRX0qGYPcVJr0FkeKsgy8B3eb3yqb0XsgpJlpTmMr2Y2mkWExyyDnmzMDfWtsD0D8BMkCxixCJ
26FFI24+MRG4f6OO0LZo/s+L0TO7pp/PBKplBL2LkL2ClnEwHBGFGiEjIikcr6ai6UrMxJm8+xfh
P53ZRvo0RoCI06Tv+9qJqvPYGLrrSqBdLu3xbjpsUxdzv6dLOpiQMFeEy6ULtzn3fb2QnhnvYDKE
AWlEqhIsJU/DFi6/N7hoyxKruzBXhQkxEza4/kcoEJivZQMJ4aFBa+HF5Yayq1+2c+vtAWcFX9re
mmVqqqXWIhUn4VuqwLIeYfYkvQrO18tRG1p8+SEqmNPxoBUNNmkFS4tuicKetnWqH4O46+oxLRxn
ErroymxINbr+eveMu30Ut5vMCTih8oy9XNLYJUBYI5TeRvSfe3fC1mnbmrreALHIr9WdJ+dvRnoS
mMfaR5gyn2VO+mnEJqe0eg7jHlcbZzTfrm19J9sIHKdoRoZWFdiUr+/GFCE++ASNkY/+X3rj3+3o
GDyBNiS1Agqq4mwBEV+cvwj86IL1D5lHL5JaVSCWwvO7HaFYT5oj1eyZsndwyHS8wXpT9xfyKZYs
On/PxWHRjA0/jWiySdHy/XpSRa5cjzvau2pH6WCH4nhYY3ruIJTfMrMq2T4bFdTqK3XEInaSe4CB
oTf3cKErVD9QZyoYesGBetMmKgW/Q3KeP3iCnpzeD07KId/fil093eFVQ1Km30qn38XXjJ2DWBxw
QI23wirah/8iQI1/CxjvL1qTfluk1IYyAgQKozI9ZXNnNxRxnh2spGsGu2OIkXUbkT5Bix66bLK2
T+04l4LQuDYZeVanNPpxfatFERzWXwoGwxmtS4YBsKsWBQ4fPDB2izE7ckbtg5fZuBPPTQ2azsve
zuYUmZpxxyHEN6pjg4cT73giDEDD+6zpCkct0ZxuI3T2SMnEZUfMjfWAuiTDUue6gESK+CJweEhN
IGndjG+4Wbs+wM0fCOx7RFXlulmdeXiXcbJGAlORUi6xe6SCka0yOA6nUuV90xs58BPBjFZWIQUI
hOIa+WQ+l84swIB4vmuVrHNIR8Ptt3Y5giU1wyEZN0mjFDAujru8OR+VUQOtrVjRsY4LrrCXt0Pt
HQKQAoH9wsuvWNuEk9z3bcb6nKQdjr8EfDu/eAlXrEdvumH7eDvw+6XxETGwYjFNNZIw5INIh6Fa
ITxxjcLYs5ybhVjP7zF+f9270kSlIIFdJCV/s/GfRtXPp6S/57JJAmiZfiZwGUCGsV5VnL63Pjsv
D5SlcicGmg/vky9o3oebA2LqCZqv0Cwpy/Z4dwZDaaYctJf82XdWhKYXhMH8zU0CDt6LCb90msoM
RVMdqjNWUXsU6t/JGW7ltqhE7ESPrEUXg50xN1umfqiqHOsVOz7sZbYd+Y1TC4MCrj0uOYBlHraD
m7ghqxhk/pnBe6IHKLzLF4fs0yDb4F2CMU79jA3hm1CV0P5xmn8igPLHFv/oxUo0lYqfWtmJb79U
EjCp9rCusZLw81FNFboEInP/2PL0LxVO2r6ryQOlp4UGd6gPpFw7HWKB4nbEU/s/nM4R0xKjH5b4
Tl30vuY+xDiBIVr0MXRVObQa7URDZtYd8zakIRVMmTpRk+r3YiwonWxd5BreF/+r+bmGRqGs16tY
++yylrdgeRb7FjMBWF48iYrOhhYGQ7izKqb/179fZM6OJPsLLk2nI3c5c5ql80A/+F9pym9G/yWx
5+mFezjfa7V6iH5OQPcEpfSLLjHqL7aG4yKXzR0TIqYVWLDUc402ZhiFrmhRXmJXzd2K6NoiL9bC
KpnMPDJZH5gmvkAVITRrCptlCnYjJiCyQfRsVnuKyjHU+V0EzEJLETd5s2A3+ST6bJn6QWX2F/YR
9IyjyvrPD0xbOPesJ1q6pulgNqUn+scujjhV4vWgNyW3IGGnYS3e+qXj+ooRUitLFyt54xciM4qa
3qDyjsdwYoL7REnoUM0RTSQmLHl1wN6XBR1wEi2pJWrjTD4/SobxspxaB55GL6ptJnYKakBRIF16
6T2ngln//5nbgj5bDQQ0GMX5nC7pRMLZTvPOL3UfSXnbAu7+didyIWGVMgu/+Kux/w0ToQO3bWHE
bf/eD9KDyQ5uW9Sa/s5WJBAML9gmV190oBeuOnMjJH/mL2PsyViE5cf3QOho+RnlkKEVGGd+xDy6
fz2AHOIFUixxhZWrh3jKXkKojuaA4T+YDz8U11zLw7ZvUziWdaNbUyxeE6w4QjIbFWeIxN87erYE
gauOBr70tMnhpbX9Hi7uvbfboaA6difz5eAtE62p0V+Z5ihpoO0YNiKkd3VlqNRYw8rAvP6rRJUe
kCJQRKJR3vKETnoV9je7YiJBU7F0X45QwgUTZw5aQ/rV66acrPM82oM7GX6sKfXw2e+qSQbdxBZH
q6k28V+rc6Ng0CYTZty7ZgxDmFjxhwQJGcN01Ot3uQbqpG78JGpSkX96T9bmI7awIABoxdmOtYPi
9opF1rh946DFHgJbv4Uq5K4zINcR3LlZHjBlfgCkqN79DP/wRl19GAGbzr1i9QmfSHKyCn6Zex27
YjUi6IsYN/uaaFRNN6Ksr3raZq0pIp0V5aH7/Us+TbLQ6vGYNSAtKuX1t4IDgsNEN6XS0X3ybeVM
HJlKUdQqxPdnNTWP6CVpPSZKUe1nvy/DhoRDIRoWiuCy13a8BtG2cwgkBI7J2hGn33tkSPzYVQvQ
b72YyL2nzUXeNTHIEfoFYUW2ZBZpt6GwqV96pfBai4Zda5W4O1OUuUnXEq3x9frV5Mdj0aCUxJKo
jq4DgQNiul1b400ca+nFoM2IN39e2r+h+H4CzdtaBJwHaWkg+gkwBJNoat1UFDxSIKgCAJKgBTj1
Ct4gSpnsFaUHQCrDoIyiYf1ZrPQpMOf8WwJ3zwtO1IR9POXe5J6otWGJjXC10mb0w/YIsNBk+Yw7
GQ0s3pbffqq6zKTWNbPOzjlE64JUte911CYIs9GxrP6gaivc+0zbLSWY8VbTvuNL1gZgrkIq7eIC
PYyXEiqqiRfICCvqxmud3joMRLkl60MSITjPB2+0hBdvQ1FAZpo4sRjNgSzQUYrx+di2SDzYQkRc
Jyo0uNZcQjacM2942+9jsxAoyLdjro9WQl3hnOY7Shxcel1pV/xcgMNAFbAoJPmjqamZQmXqoqH+
075ORPokZyM9J1GF8xmqpNoHmZaWAvFU/xwt4Ks4/1zl+jSVoXDbVW59g+6CBNYukOx6TX8r9m5l
qKpcG6JdOLIaEnJcEsgtJSq4HVDODYAXlNxF6zjdML6pBImU+sev+AsM5iEusS1zKJBXQyaXizkn
Xx9nY15Md2vrP+cnzdA5SBANODEUImJh2Le8oqsjkQfFeBpim7TvuJpWrrd8hknSAD3QC2AFmrjY
Y7ka9kCXGPyjY3pgwafIapN4ffg6uI4mcXWsibhxNMpCZtM/E703QTPH45ZTwrfUBfm+ab2duM1h
ErQtHyLmABqJuBNQx7f3Ph3RIjwx0sakIfeUSdjvCrRadVRJL9JmOzpyiljXfpH0YJs95G+Je2tM
fRBwiLpphGH4GxPSoJezTSO2UwWtS+HDTmVhFook/OFPmsOe9PXGvnXfGCV04/N6I2qXcgmidP89
Cl38EsZxfJgXc1E0pw5xVAWKHPjuL46KN3efPvWL6umW9eal/3tZO3JZmuTGijTJEN6S5Ie0Hwdj
W2dsPwtK2p9Cs3IcX6inn3H+PppWoFcam7ZqlZrWx0Ci/hKLFZu35Nju5j9d9cPXxkKKj4m0JDxq
hDpumXkIGX8x22Q2jqHJAJTTsI9iSmLdquxOYICpWYMCgFZTiTKRBNHxxg588vBjajhR8nAt2cy6
/k0CxNtrumOVK/9QRjdp+flqI+iyyY7/NYXyfGwpWYwbvqoSRO139dTRqeFIrsjI3LnFxkaiyHNq
8AXgRkeuUxfU76Oz2iLccf+HkfqfEywWZMIY3UGTM2AJazOIaCGSRlR5Gpt72tdMdIVFAXYA/1sA
g8AQ5PYHSTcwLUXganoNSSuheOkSb9LHVWbGSDI+Nor4D8SplMPwwszhwNA7bvUea64bZekqzRIz
IZzFQ1qepEdMHIUmXAHE+4tNa6KCPrwBKQIoDurDB7GHWrAP7pNfEKbx/2YrdnOIMDmGx2r3q4NL
ZryB0oySRAG8qhTJV1PS4sNtFVJUxXtgr1rKwnJT0hftIw5BNb79OFKYkrKv5ApnPvbud9tOw6BQ
kG5SXGJgMeVLvTDJ8hi5yMHqmjJRADZoDt67+rCfKW+Cht/GiAqO6avgEn2wVpOwua36zTZpHPOr
Kp3mjf5F6Rw6QZGZIZoBZTHH2wF+TVhMfXpM86XADDxAJbRCh/bwJ5rkhpODSHyNoEmvj5foPAxs
oFi9XEBwnYhYkdKbCM0Ire6srdXux0fBAIDLTuAHAQFJtBd5Hkd63hJJRudTBKuhffVoRaAFwE7J
Ast9u2KXtJhjdHgkmPXTNhEAnO/BZdRxuDTtQHc3eYUrDd4XS70Hq8nsxolx7VhTZzSSDgHM9gzN
LLlWPU/j5cX00wg0JO3Hv1JCpNnYZ5MtqimLinCYteNeDKbud4KHf+amYuzL7Wv9nCdGVF6z2AbO
2ZVVKONsl7/6nzbPJe+NLwWgmyGscC97VB428V7DvmrKybbrN2vtJ3vji8Em92zjE2+WbeVJtRe3
RX4KB3BsKSOjaCpF1T1geVozIt93X0hsgBNVXmDo6tQK94Y3HCLrNLcXA5A5Kgao+cD9ZIbppneQ
jqby6CuDnWTw/KM46EF/SsABqh5PORpULdeBfiBgcfP3M1lXUAdm/gOKWbOiMatOcl512mZ2B9un
fpz3zHE9yn/FGPzWOlANMo5L+hMUGRESHLV/W0ZcRhzrlh9ASAjzlJNezE0iFxdiaB4R/k9xFYxB
ZxRQ9dKrLB7fWLe2FDhRvFMxlUEoFl6RG+wTxkqmlw89TZ04VMcOSkOU4/Gh+87D4L3dO04BchxD
WvBvWCn1TBIZXCg9VFQ0Y5jhz/4adCZ6y2trqDNvwGhvVZ7lSoXnMJy71diqArULJkyiuBBwUyRe
MgjdYYnfdGB6RkiLc47YebYmQaERduxURH4g1zUnUHqOFGudniqAz4UWwkEVABzKwBAKg+Tiupn6
6fPuxSLy+x7MWW7Ww/PZYrV40FS/vjoNcpHuDUBWw+z4Oi+95/2TcrmyFUWPSafz0nq2ApdhlXaA
z6zs+vJauSY0uWVOca6HpnxsIDNS6Vg6YWn5B6+HQYSyrwU670HlP0PZeLwv2lkS1A8n06HFutc0
Np5wh25dSbgi8rQhoinx92bmx5WRdcfPldY13asRZGVncLTk59N891F2AX51GZ7CZ/XK++DiNkSz
MC93xDGKy9hsjjtFOgRGstu4QGymAtLBqni5ikAHBIl2dmhQBO/W7j0+tzqghClJ+edVq0pbB2QO
sTKtWYD8hRxNMcKBhvLw+drU/rKrwBp26a1b1Kef62LXLjwoW8fR07rrXFGyTE74xDyP4lXC/Lbo
GFD+BRjrmGbRk+i2XuE6oFM4yc83uHJ/OhECbvuT9uu9LgdntN1NSm1N1oA7Dt3p6zYvYyEXMow1
dK38/B1v9HGUy5qWn4tzsHOW3IcnsVoFDo1y8T/18pljuWqO50gJZTRUdgziZAfeeHKmzKiOv1sS
sZC/8nOpASB/LLtqFjE4hdQ10XWSTS1MH+xrcOszAN79N8Tpu0tfCe41q7ZPi0zutyZONxTH5Qcl
8y9Th95MJgynbfnOvrDL3u9Ofj3M/YsQlnVlHyd4WDjLQBCe7QoJvafbTZ854w5rj4p1qEErpXSy
y6gEpt4gkQNTYrThNNv+KGyyoaO07D2dh+uLKklEeiZ1f3Oy9/rm730ZC87rgUUmWzfDHJneG5+F
ksyxwlQXXnHzCfik8zWt67A0bKofh40Zx6DBXcjawByYo7so8oYkgyFVYRQ8HNU5Tx8snIg/coLl
YIiqWHsx+Gk/yw/SQO84/7axGO44P+9s/jtbN1viER8K+AU7YsgKqVjXugX2lFXJFIS6qHqEXY5V
f+lfYUFraYJ8Mm7Ewm37P120l0vjrWTj32HFGDmraQwy1FEBDO/c1sJTYsFvpsFZOLxdHssGG3aK
VSBOZcdMJB4eFjWE5U/KpVv/sZU/oOSfw6TiSQijoJRgsgKuD9oH0U8CDsF9x3Tf7/qp0L0ONAeV
C2ifaVcGX8GBm04Pr1YeNDYQ/OTaexr3CKMWIjcW9i2v7TsNXEvh/ALr48wZ56vzC8l13NjnYoJ8
1NOZpm2xb4JbGJxq/THKGFpE3111Zgvjf/IksTeWl0weRMP5R98cgMujvC5ny/eYwJOQ2ihnOcQT
RFFwJ7999HKYeWGVpsA+NOTvDt74NPNsnK3IUmY7AGyF1+UHHmm3PymbiH8DwlfiupeTq1NYa3rY
/pNHJNQkOTeOY8iKxWtZnFwrfEH79sdtBKkpBiSVZLgirT2QzjK4Ki8LQK3+azPXBaZOfRlhAVe5
NI+/0xrwgn5RMAm3s3tTXlQD3tEUz0PQe/5HSDXwtzSc4RHIsoWD1t2M/c3V+gcJrwfkIjrYZl4K
AwwIIhz8oZ2yEhtxVEmyQ6LuQMAtknWgMCCY8zT6hbTYgh9u8WgLwWHm3gK9g1AYkiw9wBzvsqbq
aFMK42wRFRUJPXiVeUU8wwdLjXANAWzmqDzShzvApSabvpeqVrS0u0CVTwsFMsINKbWhDbDtdPUA
EgNnmxRz3iH93WnZ8v68jlrEkHfw0+krP08PFiIltEp5UoaL4iGlz5b5nR6dAoP5l6Kfe6Hn3j/2
NKLL9A64awc/DWyYGFpjZx2w/GkSPQ1nkB4fJfJhBagn5VYKK3l46B/WjQFCGm36BdTTiBRx/tsr
gInzMfsZwAA0XXNHMUGYBecWURBt/1csKz3o4QMpalhrav/M6XUbyGPSyQKh7MBvqnWVyt1cZqur
7eS0yJRE6JLToTf1IF7Npdt1cEN0kcJBOVCbHFZyWOit3Bry540EZjvfeXtQ4IvvGk3AlG/jV9Y4
sDNXSdlwF4MwZz12T6xclMlCoFupaT6FhqakPzJL7vLa62bN2orSe12UhQ52FhWzuPJ4lGUTV6pu
/0nYvmTGFCYvlvb4bnax9+ZtsmCC4vUjizW0izguGEA9gFNStTgm3Wrc/SVgo2m1ownr4OJO4fwA
Xz3lTqt0k6PjexSixhrcaid6r+msXIu+ANtYvpf7sfdQw+42wrNZGyezEkUsMbaTDcwM5TbG74XZ
9gI5LTNn4lr/aaVta7UTI0JcJapnYgxZ//INSCXedJMyIS34pHLMK8VvA6UYlue/cgijSZEAOwl6
y/31Yr6NLPAVyPNXfEFxHn/CmpIXuUQMKMzS0YtlB5nk6ZgEBbDnF7lh3+i+MUwjki4wt975mHqZ
nfO7fFiqCKzS9BpyzexgNUebvXJtUubFFKW0jMXvgo65cLLle3ktIcAtrG/Vb9sNaXgWjGNnVQ/u
DQ1ilhRIBf7ZG7Qpy0Qwk1WNVo1ohybt4uqK7ccq3uA8jfnVYUFEjY2jpybh1MILtGRKis3KJUfD
PRs+zF1qtcm/nSXYbqiah480243pC+GxDnuxHVVfEcGifR73Z6inNKQjqPBdHBI8zMYk2k4qAnKi
tiekvnYoYV50KRM9XeY46DS8EO0xablIwjBTR27YGdOh9RemUsgCLnMId6pDP4luJAibJQRpbPS9
FzTSdzYrVP7vEzeDZSJtHyLj3LPOsBNmh4aTPtOKMzcipTYkptZbMqqDKuvAEX2KxCGe1k9iQ8zr
2cu5ZJyw/vSuK1DTatHYkxTEDfnDqSSlgoQBcnRIdoE5AWwa/qBnuLyjIN0DhZ67cqQy9rc7/5Hg
WuSnIs8xjnz/AnCDp4kH19GlXtq4QpkdxZ0bXF4c7ZG29hPKekgprrisrfl8pPFA1jrfJ4PdNzE7
dMJidXhjZ/b874eUe0ziV6jrstPF4twDRpWUpWxPVqFGBkv8JZ4qzicLltuGHBU9wcVbNEyL4QgE
F9VyTfDWMYkzeYAfT2BqgeEVuPRfWipDFzXEBInK7VebiuI5oTlDYeXpX1IHbwt8GXsL1KbLvgJd
n8UGw/Xs1P90D8Yn+TyRbj27zQuDPjmQfA1tkJble18EwVIfHnDGQh0aDYeEOZtHPXo+ST3BFw+m
zQTGa4gRCEK5dZXQE9V775Z2JFalIn1+a6NtmdWXieJUI/QxrC0lyWZFLM5Jmn1mh4pCWsmLAbAB
1PvJsS8ZULEFYxe/yRrrILiuR+blQNvJiVVOD9il9HTBRE8YiTYa353MloE0V+ZCCTgroXoW8wVQ
FlrgPAMBx3XHkO/FQ/pmgUo/N8vOdFz4bPIWPTKvxEtkPxijudwwhJHr99uqoWs6m8qPsAtgnUAl
xlriXNbS+HroEvsZ4FacxQkVTxPik4oXnvT00tBNvYyc1EAgP5MUatDcY2DoTY0B+EfkeA7wFGG4
nMyJcMxNYyhEbAU19DLHu2AOdXVav1ZCP74FntmEH+QnvUFK7LxK6AiybciGNRvcbgFcN8OiQ1+/
DRuPWWZ4ocKxZqYzwIjRhFh+dJbYKo7zt0XN/8DbACkzB3FffR02MalWZ8E8aM04tfhlDn6ntGQz
ezJGo734fma12ss7bCvwz9Kz8pGjLddu2TGoKuH97QbpPBjmORf2AZ9LxNhNUX6j1aOj75jv7XOm
I3clW8FRO34oWolE5PQkOq4q8E3/UpfKndfYVgHIyneAlT6FAHGnw+35zfl3+E6y+NOiYrwd0hKV
3Oqwn4Sm3v7+bm9/a6xIDoe+44r/fQkJBJDIwmu2zN1W59q6j6ur+u8sdtcviSQpkTWVYwhLNtbP
6y/UrmPsTxI050p0RZ+im+PeHVJ8q6nxZAZUApFl1PDgcETJ1tk3A8TwZ7f+eT6bRuxlG0tdsivD
Ex1mT17ks7kIJMWBfQUrht++6JHNhZEvseXbflQtm8dW3vFS1O5gy7B8Rk3GObPo5TPzh7n+5lq/
ZKPlrV4ms+mB9ZB/DkxtJCQaucYY42paqg+kZ/pop35gR4iEk4/vucgV4wbrMvbe/JNlXFciSV47
ucC7JumOhlbJ0zxUl1vTMyV58eK5AGanz/t7/avkamRFQf+k/RNnX27JR4Dch4JspDJiE+gkx7xQ
Uf1Fd2+vGU4BT003rnxL1mRirS+PZpgHthh5O71mjb1NKbuOh9mJS0+NsPC1elu6a2I5tn5jIKug
BabBYy266apZDe4N4QETPnl/+oDbtQIcwyQzOfbrX3wMtGZgwmrL0erAmrwjA35mfxGvCN/r5fFo
6ZUVKz7loPvmiXZj5RkOkLW01c8oW8mD9kLEGxbXMximcWyk6DxMSFKaB2RJyeQFxUQZLeLYeCQI
JguUgY1z45OyyomSb7+7ryvRM9syLgjo99J0bXhAh0WU8MJuihhVipY6o63ZWE7BV+t6WokIwOQl
Xh4sC50vzRjSYp9+OwqfLhJ+9vKv/a6Ietj6FU8PRry8bfLwzYFIebW1wYoYa/xS8XUCWQ4Hdruj
HK+t58kriGa05b2Pmwk+OYrYiC7b2sb1N0P69hWjInkzYqcU9ilEJE4v1VtAnKcLr4V9qDAuL+2p
csoJM2DtpUfWgU7tKvWHKoJQaxqFzonrwFzWIxEgey2mOJ9KQSIaS3TT1UdNUPKbqxBRbG6FxTp6
I4vdwJwG9JUkDNakE2GzcSMntRqzKWEmMBSrtzpIiFrP5qcTQ8Tr8cB36SDuunVRSumkj/Y4vbkI
wLlBf5VIl/QzQlj7nbEM1xwoxCsGufK+eF2vy/IdiFA/iAC2LZD0cUtFt+wqAAPSQESF83ZCmlFA
/KiNcJig6HkovffkYU4iLIYmC3ZHNR4J9vrWwHneJzEF24ZzDhlszOn87bxfb2to3bHJdkFkBEHh
va4JxnPMWPZlJYWK0nUT83Smjx0Sv5quqYXbUydACWyZzs99K+Zu+PIFv2UZDcTCTezSQm1RPsYn
EPegVctMz/k6vc6YmlXh76xHNKx3/JXmaFEb2HAPjkHfQxJJOAYEIh1/j5s1SC70Pen0cd2U5AGr
lFU6WPAXVd9r8Ez7XIeik4g39UMUvINYhc4A6UokjQnecGarNVbpwL1gRN+ZZLtrDNlGRt98uN6F
B6gmGY73k7NnBbyXVLuBi4+04TUANSnfYDsO65irr/ha8WUymXvYwUQMe6S2/K6iES+t7t5NqFfg
k1y5Q9I1XfVW6ucEHamS4IGR518bPgYNtGl8Nd/yZY+9D72cEQlwH2zNCliA/UyLRAEtYCms4BXy
tlzNb1A5gXpMkQOLaUv8N60m93uNemmYeegwRBEqxr1CCzlBaCR/cvNQxEz2/peQCQ0wbdQ1JE9p
jpyxxMqr3TXCgYz2IjXX34t+kQCiTBZmQ+D0I52531Z1gFyb950CEg1wb2rTkJ8htzqMCDz6/2lZ
MKucaCV0VA5mHDI8k8X6fQFgXXXvwPUQD/Vhv+6OU325ZiTtL8h9JNE80C33X7zAw9/VeK5V9PXX
d4BqGSMgSZXf0dVv9kaqCgH2lDAdfcdD01Uds1sLintWnmpveF170S02QyZLpsCRNxcLvvv4uGwA
ACQlh3B0nlMIeVYUpJTQPKvB3+yU4ZnLSA8muiuxpfoWk9uDne1HwczlZ1oxGa/V11bPyjM3Sy80
05HjyUu0/I7v5S+VQTTJj5NM/civhlCPILz6KVVfjC8EM1aC0mjrN21JVmXvIupv6fqX48FuAr9G
GCY9wZRRKjRFzLtxgiY0ImqpGq7EoaJ3Wd/1L1f198EVmMUZvKRoZIS7lUKcxiDBGARublooVasq
Nr6jiK6vq3botvyZ5W6GZR54dziT4fmEmJ2g8nNjx4JdeH9znAfTyyRDIBbPmcOKDZQozzWD24dn
5+jst5uRa/Xl8zFOZRprhx4P4el1u363kD4aBXxZUssgH3pMduLmF89tGlv5AOa4JsOAWyRgVcKC
pKFz5B1wkXYIeSMpltt4bSQWhslaQiMqPlIQ8PfW/G9Zr0JlxgTbQy6Hxhi3K01VfYQiPm87CnLk
JqmV+8TLIdx/M6kAZhtJBzmOnBQCaA0VSB/KVpu/OvhXwB9rBYzbiKE44KZkXwN/JKku67nAT9wl
6JzcgqaRpyq9FBgg4tCC5SFCQgIcE7VVUbkTgs6aKNLF084sTIZD4sNO32pvrakezX4IlGGPKdKG
zCERglzSrVmSHWXGhVvhgkOybvVTVb3z2DfIWG9iq84dq6GdlROD4VXdC8098YNVsmPcXysNDXFr
ZO6htg/FM/J+WifQW/JXpVU3scjJKXW8gvXL0/HUa2+oh8BVvTNRq5tKSMdg1J7wUkMHE9NQO8hd
/6vt7ActLtHqzzF8JbfLumagN55gfc6HGUgUDt8U4CZGztT7Dozlyp8Ya+dhY4gTGMLxdyGz3de6
Nh7XejpQVb+ieXbDMaQvr+g7L8gMtSkwd7UEEMM6Wq3nf++JHf95BlCkFksZQfdw6cO9c45kgv5V
sozLs/JAXHgbW83EpTj4uZxb+oD4RPJ1bN1TDJPNJWEs6DpBFkCaVcXBc60+95mXzCXXFoPaQK2C
ASPA04Z21cxey32tgCYkads7HlEFIRajINereaVMWSbuRG7n9FMewhx3EYxz8dxz7lGfnEP3/qUs
QKNX0DkmjoBc1E2XmT9w95rem7z/x3ginuthfss8hMEWAkRDbbxVcl2DGh1Xgo7QQZrcJ4R71nNx
5WhlL8eDCLGU64Fi0dAhGC/09gf1pxwr7LezZRgwsgCyXCKkwwKbD0SHrVhDNfx2QbOYs7DGp8PU
zqmuGiJ0JRuNyE3qX8GFyJapGw+NJw8aRZnBgnrlaRuzu8kDF/KVWq76E9dYl2C8sQbRnfTbJMpr
DA2l7R39TK8rFHI5Ja4iBqStuaqQghc4w2/a/mdGIMKSM59tP92vp8W/oAQmp5+M2Cf0wzeY9puc
D7t4DgagEbjGEt0OfluAkEp0KJE+tWrwdxXDVswyUKhqMIpbbnoSn0jpGy1BJF4FG1qdvvxv6/3O
pG/01AtkpDmjDOEeU1VnlTOUDFHCIYBfF42hmgOTzU2K8DeJDm9VEATshZz753I1y7glTAobn7xF
XwnphfpKVE+V1lQkTMX8YjrDCe4K36qT8Mx98FzWav2XtidBC4sNvjyhd7NSAwLu+AQZkRK6MKDF
2+qg7VfPFYQNfYmqf20Y8g5uHAr8N0D4LWzY1plOBL7w1BvHUPDT21/8ZVgM81TBfX9ESK+9+SEM
M+dHEdAcL88O4p4RU33b6ILdv2WnO22qjD8pwxw+6vJkBR/F4nYciJorDvdkcG0BNL1PT5hvktLk
+pEGBOgWrfireHGDf2pHKtpQNjfuM1ijwtJExSvnBYjPtzhU6ikc6ATB2yN7sSZ7wF4OngaoSJRn
ndaEZt2Qb6RWpO8tdiKg1pDhexvQn0decgfTIwwMu1iioFMrqGdUntBN6reM1ICadv5g9omSLTMa
PBYEcvIVn2rBEHRd9+obLCHDmJ/KLfv6QFudUCMuiOAjbHtZrFzN8htoN17gU8JGmSPNPmES55bH
Ee5zCD4WMOYJNti7i2cErlLLaM90haChppj5DNwbJ7K4LXioEPQQ3NvDoN95FEdMTUf6PIeHzDFh
e9+Ye1ErsOPDFIJvRl9sIKFimmGzHwqowkdJnYyEYaWOj0FyQpXW62is6ob8XiNg6okUmyUhRUg0
T9eC0SJa1EYFQzQelVJfcABdCAQXZnO6o+50XnUw8thGn1OKH1s72gmYJklNyjrwO77d+IzVYm8F
cDX5xV7s2iZsc7K4fQKi/jwTsonTvEaKNkubgAkIMrF9tHV8TsaiInPhfh+9aE1RWzYU0nAFlYak
1eSzVeskH6WZbaDOdROL/neY8/yEyH+Ir0sAx+hSqhYS7LeFwUTMnw3anhYzWTBuIHNkVnRb6mTI
LUiaIysaNgipijB677y+gdoa+4u45o7Dqq15mbGboUoyfkNjjviibbOA3UaIi9E4oY2Za3UF0rx7
Ji24XNqeZhKUDqGKXLfvWvLb0lPVvLQRZCnV+S92fGv7eRLNig6nw5YWeib4gLNHZ4uc3LfBp7eL
RdhF/uO7c4wggkddgswtOecq0nW34yv4ZFcdvgV6PFC7e9eGgugU+0cmyGo974Wbe7NOFj5Z8Ly1
WqJnrDEsmAXL6isBXniNau+PGD8bSL+TXZxTaG2WXFvUIYBamhMPhgOGgKrUx9HGOTX5lZlCo5vY
+ORa+Cm+GQ5PxPryqHDSXTCnsnClpeprqXbl31yHMGF4Y3bzZkZm8iU88/2iQ67+2a1JYyUG2I+W
LLdu8Bj6R1VRDXlwTUvPcGyRy271qzTJEoR91uD9efFACXZv5L+zVu8dxtszMpliK5PY/2kGj7qU
V3KMQPfieX6WFA3J1HkjtMDSL1aAJAKQGypSKb1rxzZZStFooKeyEmUmCcd8WIXbzWQuE18uyvly
eT00u7JxqGhUKkyoa6k1EQEoGYnt1fXoNRjS2wPEhUvoMUpRy1zUi31xoz5aNHfvfjfPLI1Z6ClN
GnOr7mS8ZMj9KG+Z4RAamAXRcfiMv/iaDoE154hAn37keaTYf9fg/u564S5keI1Ris+CLnbdmpAi
41JBV30JyrCylQKx1CmNxwer2ZP0NIChRDYIDXpIA5kOxkjLML3r4a1I1fkNkK2RVg3ZPD9Ybe18
RqzSm2iuSW6a1L7/cz85im/spCVnWtpby8HF4tIYDVl7gktE0+YNGGzT0/RZVj9GOkgOC0h3WTkw
R/0A3QhHAOSDKPDfdnU+ldGTAcghZSVxrfdevgRal/ey1PSNJXk+IU8mKt4o4UNEwUPRhQ3pvGps
kzSPMDnRZ1de90PlSURx2Hzw0sv0NCgJHceAXxqkqYqMrZkLQtM4hpdNsiOAbfe+ftNJBmAYq9cd
mEuo226P9z1FB9iC7IymGa7fzXZ87vwlsvvGrcYjmwdKbXHlXVhxFHinqc0plfDdzv3SKFiQwYpL
+AnWYe9XmTKgkGk4uqOkjCpc6YIv7swqzZ106BbNUe6PeS3tdLYyJTZb+D0cnY9np/d3tQyKRdPn
JwOf67NirKEklOKEOn/j/nCz6eueCSos0GYt01oETAFEeu9La4CihQ+imlUmYqcHuVxtohPXEhBG
7XnD+g1dxhf+3oq/kMihgyVYXfSLBZ6z1zZnn6IvFv0ubXh6ZrsjZYymyd3Z9dP912afXAOCUHq4
JSCaZdDvYpNkT4pKDKCrwWqITz3MWlodkkLCsi4deMx6vYvRgPUxQhuEQVvd/KfpNWVTb0Htg7H5
9vl+XXnXDnb7fwtsxf508iOcJ3u29R24kVV1RqrhBVVXWBNgGJPjh0JRlqibIWOdrsSy7CZmi9jN
MmCvQOW+BUXjIeSiR1SqRFfWX5ko9T/AqyED0LurKLt/nxnOtM4Vrtms0+CJ3BOdQFa7vOH8llqH
p4pWU3C2BaCI8PrJEg9HWHe2ObLsDEAHruvzUtdm15NAgO0P0+6ThsOI1OPA7G7eNsfUMEmHk013
jdIhnfn7m4cYkmVQelGzo60k+eVBRJwQXf0JwKqhpo2li1sKVouajAL7feqDE63pNuNJ/Tti7Inj
TJxwhUSoZPpZRdurSsidgTRkvbqj5vDbq3jfVagCarNypJsvYfofFUj7vaTfsPTZ6M3AxWgpQl/h
SRysLUk5vyqhlwPZM+eJm7eLQZiVjs0V9mt7zhPKKXlyb5ZwWt8UJjtE/STuWtAU7hZLSh1uyiCE
5nqmQrL/Uwoq6MsGxEtCK+Xv7Dcfy/koFYiX4tsFjgBfWzqjyAuaxQ/lAIeYg6MMNjVymSXtybMm
wGfDDtU0pVB3vBlwhMrjy490tp4XwzW02G2aAPOdu6HkALqbOQEw2Sben1oneMeJDMiJK4arGG/l
gJS3rKwp1v1ew/Y13tDSgFIqkMKD4by3ldzk8+W9sudiE2HHpDHx5z5JlSpoNxp4FgZ7MCG6KN4i
HrJ2FnnyVH1i3Ox8xcDBUkmSEwb7v7XkAsB5bq4CSS0hYAfy2WpW/pb90qehNGhzwII9Z/hUNTOK
xQY6vVRHlUQn7kDNyjokb/KRy6mbDcv+lkcd0PgZbUkdZtk7Dat3GbzJz/i9e4Qt0UN6v9vSjiBp
4Pqd1JCD18yUy5va5fcxcVP+iFG6kNeQf+vYpBSRJwNjtXhzVQcS1DVfhhXEMzFDkAse/q//RlCZ
wkAUcQ8LpzxdXf/uQzx+BmG3wFkQNd4SdnVw+eWRJ9f9vkRpQDypZ1MIfOWpkPjksJS8wtcCK7tT
5bjXJTgXbjtLsmsSHr7KNGjN3Mio9JAcHAMxNvTaP7dOLOxHLCc3YioDSg1Js2ElqLvzOgcqG4nC
TdUn1LOKB7+lBTbCzoTm9a/cAczvc2CIotkRENZc56CUrdyTA3qNvLXCkufZNmaIXBp0olAYMuWR
Z/jZA3ARfC5uo+/zbr5XMPXqhyZ2UKY0YSh4F+iEVGNvkLVZrZB/iS1oNAX3jDslJde4efmd9ca9
6nrV4k/1356G7AHo4cMFlrXuFO2dqoAvHy/SG1XDuHS/9ZtL5P7aRg3iuEYW6KsRzLe1p67pRsMZ
TJDreSbRIRb6gwhW6hyF3XEptYIUJP01QiEFle/ugHgmskyga7tqxo4R7GZ6BgHAuasW/EMhID7a
lcGlzS61SCS4sv+dPtDjxiY/Pzmbns9is6LceXwI+X0KIMafXcSm/A89lRrKNE8GDALE01SQN2wh
wD4xK0u6xkpaR8Aqm5DYV6FSteDWlvGc8t5+93Z4c0Bpu3yOX0HUS6ETO8nCDgeu+p7dULnz3gsD
FD893KVnzr3sXbvdpcVmoNHzCt1FeRtuONLX99BXTUojk/KvT1fXcYtF/7tEO/fCxhjyehv0CDh4
XRQu159PYAiDTIn4wXofMp5oP1icMJ5hZnf/EZjfq9V0NeMMR4ZKLpMyHGDKsTGIOfNJ0cH9uFaE
PyCWyJHKWiM43m7yc9vOBNF7A8PSZSXdB5QKueI4SCHztN7MFwn9/eAjFcswD0gd+5z/qko/1ZAM
yLIg9KKWf3qkRieTCHrr/+m1GyvPHXRu97qTkG9qFNX+bHhVkYIxIpZzs9cxYIbY3Vdn5C19gLrc
V9LiAM+oouPPcGLG5Ug99tzf30aWSGbl74soBcDigV38PlNS1YrhXVX0Y0IDnB7pbmUT7nWumvm0
SaNxJvXZd5NzNGmXhdV6BtB0kUayiTeawQA7igifw+HO384HqS9VgjTPoWwlfu5jCc5i3DvP8egw
tK4V/SERR7PvjQksQRw2+17pDPrCpqIv1EF5ROYvGf7Qd9ni4Le4NyYo5ztKfyzAzPUC/cYQWWJv
KaALmX+bMY6zfMXCiNEhkWVsp60l7wOjLOstBOEL8m1ud3ToIEIvVtDSqpg40ZQTW6Hl58ji5zW1
rNTtdqVjVBbVc1J93BQgtWGNq/s/unrJeQ2e8/90yUYAR7lOBlCn5kIjH69ghYBw3J0GKWELutXN
RLgzVgTQVQ/sHFeZ996a9+MJnpSFRBbJnME48Wch4bM9bN9Xs8901Z7ptFC4EYNI0Ki4sGsspnAh
gv4UBgbP0mGPVhpFMUAoE4zlATuJIcGoCYWcxukZzvLxOk3hWejie5LOxKC1Tj8B/TJdxeBXa5Nj
P9i6IMplrO1N5u/qcYeHB6vVlTKInS1TCpZiIiAhoD31NRhrvYWAcpJs9DfJfr59AMJpwv8g/5Ya
rUGaGbW/Dab1k0xJwYmTHmoBt+SNSUoEXZEqgcSAKoDU2tGH7F3nTXrGA5zdIpDO5SDsnIsmg2to
boXdaLrDk6p40iNkCQA6wtN0ksVQYkwdQO5N/pNKWHizW+8ginLKUVxjMEb/hPb158pvMonI3CW0
fKTUarGqqCOs3U+YjYzRdJ2034mEYDyt7UbCxY4mvNycIeL6w4kLuOyQcmhij3uVsozjaSSTRxh3
ASzSjglbChLeoWMU7q6UUUD3E70YBW1N/HPMPCIDVyG0jzkAZxgCBybXRAPiuWL1Ym6bm9G2hNuw
3E7VjGyUy/TDtvifZfNB/lfE3Rk7aSR6Hb7EUKgeBtSUfCcRnQLdRTTnri7BmfNmcSt24d+KSVoG
LdKU0cSlfIH7xm+NAdi7fwgmVNYZ1MaQFO63ZmVgGPQJO6uu3AwvIzz3VeVEzDzKp6nJcZaVwIpb
bxq4wc5ry9irDsF9bRD55+fOCgFA8mavsrG2ijFo7HWrdZyMsO+IUbHJiCfMSXnEvSJk0EvnCz/C
MP2C6080a59CHdf684tZ6hnVii6jBiHezA4zsCmC5t8sH+CnfNSAUhdGaDAx8xKM8ARr5L04qvPb
2i9IKFAaU8yzAWj3QcsStTErAOW7qbbaAUrNYg7Gr2Jzcmt5C+wCtDZ0uGmBrf0/e8qV0rWeAEzi
tK9ImdGN+jUqz6d0GfJcJdGWhCRU6wYsoDW5OIp0dnfoaZZIsX3l8a+bvVJ1fqjZgpwwZCoRzBhF
NHLXEQH7tCLgkyppwxPu6j6y5FD4d/bSmphC6+HCU+ZMU/xrKiBUshktc0szSiliewDye+HSwVQB
4aiZEvhnhvGSRQi2yhFhB9s6WfOdfD1akmmITTkGokEYLcyX8lAHkSC92xt/iXD2JtypmI/oWSL9
/ATzXcV1vSPsOAOPgZGXmGUuvfiKUD4qH4ADS5fnUtgXIvT6Yu7g7aoSDJ82qqzALZiFvkPZhLY+
ENaiJJbhnwKerqn/2RRXTM6sQa52pWrwIv3E9ILe4jvvMx2yEssso0uGYHy34Oaid86QK5XoX30G
P5mPAe51/M3KDmeI7nbnH/cosTAWIql+yQHQ6fwAJB8U/2wK+rvoHEwZ7pUbOVAHCCsTKhID4sUr
KasXMWwXBYOiBGIsDYme1LYUkw54luwQEttHhCeRrrP4+0swUQSUHnmOcStZujPighjjpe+SX122
xTbdbE+ZNIeYw1Njd/Dv30cVWxir8SBr25Lm5c54DPu5tWkSrdII6RDuy/q/N6oAIc7yM6nIObvE
EYnXiWMEkZxD8i9G5UpJc66nhBWBzf7/GVUmdWP5UR0iV9ASTQg0HuMb9cpITddXTfA8sFa+eclY
r1pUwYiV+KAstrmEOpGlGcJbVCQhgT9ZddCGVW93TcvydbuueUm6oHs/dlAboAEKGDRFIA9OUN//
RAn9YlpTdJoNX2C9FDaaGitgVESWZ2Nf1gd8U1b3mT2O0tR/m1kkULE3uit1p5zfOTCVOzbegiVe
CXXPdGm0/XuLlJLnh+2hxZkijBLs7MN2rHH3Ln01kj0l5hO1EpCvbkNxB6uxT6j0MchIg4RWWc4Y
95NHcPurh7MeVyXnSkMsI9dRHYtHgYWPk0H5RvAXQBt4asMDtCAgsXbUss/DX8ZlDMzitXvTbzl3
ZmoH1laY+dkGYHMN/G90c0Fao5T9kiOIAJCahR2W5CypAzCCaBP4ho9qLC9fjAjz2ISRfNAk1O+O
ZwlPp3nBGx8TXZYbMZUm4drIx+HrTIRFUAljmAohJJ2QtiSuBb3TNQHf0Q0i1L1wnRp2NIScMFZ1
Xk9GflOCm2V2WR9Pwlw1knfMr9iECrj6D89KKabaNVQXbzPfgVG+Ol8HrWhThZ4DUtapoValVHIy
tNwkRLOMjCrw2ttSf4jCA6/Lc2DGn+nM1M7rejK4mF7u293AGOsL4EBgPBgh8TGMyLPC8fDfkfKv
b9QagH6fAAnww+O+bNHsYR3bQwh3ZPltFMre3+Wk+TVG8f7KHWND1MSc489EwCCIqL18rQxbCDmL
8D0y4EKmscLDUs7AEtfcB0vQTySZR2ymr4r7k/BG9NHhIKOf1Mep6q1ZrDpdIO0RxkM78pxeye5H
V+iA2hVf4LPkVjsmsK20VxUk4iRGUwZJDzGI9rneqrgWATq6aXd4KyILxSZzoOLxp5HOGrv7pcov
buo9ZR3jJ04/g2eEjfu9VKK30mCuDzUqez+Vgsx5rTH8z49lRJwPrX5mf9eYh8b2iPC0gOd75uaQ
LEFnZuExMn6c36yNi1NhD2DCRxTlOmLHPzad1X9tpYNzlks3B4KNFLmYxZHev2Faz+EkbF1iqZPi
KN0xBYf8k5VrnkVujiDPhViEGHul4I7S16K09rS8aDYCjuNu2lXb1yEQeBQciNXrMlsAwhURaz1K
1d2U/yAJbsOwuQey7gxsNLtzIM3OKsghokcMGZUt0kq8+DF8ScgCQOSXW/lQGgnG69fP+dCa9sYr
SaiN7BgUa68ePTc2/cCxNxiw7YeSzGQedMWJSyjzViPwvedertLeq/7Lz5IFW5ZvkNiTnSApgm4D
NcYsCPO7JObWRGdjaEW5CyPIYIIDTvGX3i0QLcvOjI/Nfv3DUnmqOTbIdcg9fj4E7qS5koA9WCsv
arWPzrtrYH8VPQZd4+IUwoF+oeDF4cWXmz04zE6bPHjbQRDDkClXTUDnqPll7ucUpqA+S76tTNRt
x/4h9B9phN5GrCqjVoOAeRXFvYt4FUAQeJIWGpmEh64LLQUMkYM9IRJq4DMQ3D337J8yCO/rzF8L
KishCsGLDfakKZaerirLIxbu/TA2J/xG4NCiAZ2mBIhe67ZhHccHLsj0ICGG/or2tDiWkTxMg3js
b4/WDlAMKSLf8uOXvKB2I7FUAQpC97eTxlPtWA2JR5IDNctgU4NHdKG2Ih8RXx23UlEGyv75nWWi
1okp616Z0/gb+31s2wuQJynku/dAvoCTkJm6igaKmBXJzgpFcWS+0QvH3LzJnN3niTXDZCpVPLNf
XDMeEpvGEzHW9Iq34udEzj9aL/SoxWZAfpFqZN4gJ3xByu+pueMu76y7yPzMCfWG9u+ipxOQpE6k
rHleUMS0ZUOVKwnD86OS5jjtp5Qxlr0zaTzaiz3OphEFtPl4EZVJtG33mzv3TJuochuJzUdYpYZ0
uCvElM3/0xIA0sBtRheXGE98m4OfCwkHlwXkGpiDn6MiRHB8lbrvXpIsd1iuTRlFqWNPnvuf9AQT
IJpUM3KWZJ5eoWujONk0r2aukivhXGrFIecH1DTCNKXBPUtOrAgXnYd1+rjiDQ2H6NnRWv3sA8qm
0HTX6yl7GcrdTzXLmGAdvipGqfar+7ssxLHwAiuUIKsn+t5d8tlrbCA9kaqGJ2DQF4OGgEcn5c5s
F1j81QsNLYjgCcI7+9waNfFY8yYTfxYChAHu1NBGJjGB7YXDY1PD80iQr3naE4SixyaF9tMnjqkZ
qq186iojJouvqIgPQIEvjx+VqvOX5YGrEkDpJBdWNg40OuuOTX1Z9Lr7GEigp41S3EHPfcAqrFjW
XFFGOpOIaymxFsgm2LiFmcv8EFTynGkZxgmRGbF0nAscC/4cj3PFSaGB9GMJVucWVAVei0zZGa4J
xG6PITtlOCMlogzlEYQ0ySbTEU6foS/xJBf+l4hUSdqE0Fed8EWmHY7hzNoBfrD+kd+mf1shi6hM
HcWZTk+vCw5/DLjZ/vPjmLQXlrcFEBrcp2eR99C1pRRnfGR6+bRBJSvKIgVvEVTFAXNnrS3QITa8
LKdWX0LdqQJkHZx9YL9Bcv3dMZQeyTlKZqi7jrJLhM6k6X1mTeFeSbAX7Nuwn/LaDRoqQLLj3UA5
LZfhrJ16NaV8TgKx4W98hgrljvbEggOZI7oaR36GE0Rkw3SBmtima9qWoy8oPs8BxA+Vv2f3iw60
wRxiqrss1/D0zGosVsg9xHA7DtUg8iEEJzdbJL50/aGCvEEnGTPsUCQR2InOhWoorY121m53u8aq
WSixqiMRGe/jbIea7otVwsbgGaRgupO0uHP1uvpSR4YQei5Bb3vZXkPWIRo6Ppz0JHjBPr28JZ6B
5AGHcTTBNcXmRv2FH3bsTZxnAYhNucbXxsII4fshuMAZTHXszTRiELz0FduhHY6nA6ee/o2178xr
Mi/yccyzC+J+qGzfNdiTxS9d8HmF8qmYuNzYDbfGaj5Pz4yZrVYcJ35seAXB1IldYxzsUKPqa5ZP
zeMX6Sc9UnKR0nbCg4C0Kh2t5ugRVFUA7DOL4ko46LZ+6QPfk2CulpndkOOWmXr9WEqiA+/6jjOr
3CQS8EYGJ1+Sks3fUJN6rQ/WD9x2q4xCvYAqBClyERCOQKNs26+fWBdio+N/ne/yV5XKuyQgA3jx
b2sEZOYmvN3g4mmVyARJ8PC5+kuJgG32ZqAJ7RJvCjHqskW8XfUZisT/sOL4x/Y7Gxvja1785LfR
5uM4ac9JyvPciWd0/+B9f+wlGYUt+yfUos9xMlZssy/bkEGmG3grF8gBoq4OccRz4rCSYWIx+crP
Xgn10sUHbPIywgL5DQcKTWOkSIink3S6fyMQJNBBg1teNfH+HCwz6R/vsNHGEcTgoEvo6hq56yYc
RTKqE2czLoW9DdIG72ezHGB4Ivc6AW5MvCbDuVOLSrpW5IF6VkPZiEqj0boYf+I4yHA54zrLWUxR
nS4KIU1Lph7zZ96gacBs3Rj3eujKQHhz/0UjMEnWmn307XXVlXkgHXcJ5rbRujNDcyJ/pLSQf23E
LvZwz0+BO6sn+Xzpk7h3r6drnBqva0mXe40ExoQ3UOa/25nPaKdAHShhtUgqWTX4AVXCuh+/TRr4
3RsptKwC19qHqLTsedBHuRPGPL04lLFCrYMMGjg6fhEEdLwJB8xMDz9vWC0ZNS/RYeAU2Zhm8P4o
ya92LG4Xji+cWNUwjR86HgvhAy+KeHoxxOQihNp2Z6oNn/PBoouGK/Fbf7IWra45UvNGjT9ZtPEL
qExIwpG6hMk3xzuO1hhDUTXa1xZSSg+L1++4bP/+GmwnWmNmrcK6rrEOnxAojn7/JoU9wENB6doj
7Cx5nuRomEuu+SWNO6IbqcSqafNHbtI1hy/jkFcEeqSOBBJvNeJog9r2JY3AUOwSjIqYC2ca7SPn
PvPlaMEKBGagZJOQ2TVHhof07MKxJ3zZTs/+lj2tFQAorP2vgTqrv7P4QLHDHINaw+AadMel6xtL
CeoPGaXkQTT8zXevJcJ62Lt6gaaoKyJairOi0E+EZbo4Fl/It+vqe/FOnk4ywfMZYRJX1soQKdlg
uldyo+quGMhcjSsFpn3cUq+znQAOQP6pJH4hWNxx0sC4Yt0vPvF1NI7ePdobWTi9LmzBRMYFephZ
JGwQ9cWfwin8bIW/T2wRioqsbGbUW/h9x7NUFbnoowjYFJmTa9+J52M92y9G4B6m32yH64iZroQi
jSGLa90ksEEYbSPMBD5OQfUTDvkjYKZgS+gKUM/3IXOELUBOWn3fwUJxFF5aVOnp+wWRurgqWFD3
DJ9ws9SKybwio6rCiibgVVaeZV+PXTun8Nx7DprtvoqJI8OUID4Z00wN65nx+xPGtxAufTIpntWP
ryeQhiRBmWxkVzudaJAC/4/B0SPANyH9en63kLnxrpvJo9Sft7h2I4lfOS+EznL5ULw62iH12f+C
NM0kC/Vum/RBEblnbYd3JzONf6Nv6Zlyzm1OEJm9v+C511FvCs/Ik+n3v/QUAvDCiN6N4/OVeya3
dGDIvcxyAknacWQGwLhxDXgJxSsma0r95OpJa4VzU0qbsOvyL0sQzxWm/kJzR8/ziSnnJ8TzmInN
Uo1NE6yLgcIgx5czeJVgbSpSB8NJvHIEimpRMg4zP1A6eTd6sZPHGA5NQwxq6+Gkqwn1bmQWmONs
SdxG2Gy/ziW6v0h6T6B3Hy9r65U6CdXTsGwweyknqrk/HFtQKFVA3ViTlL1lb2uhSr1+a1u4CZNh
Q4K0KmFwtnjZ5eXaToebjGqb8euKFPnlDo6foEFjtRK3Y3gX9oX1PIAEHs7mCBgqjm3h7CWH26r6
cgJ9+Ycz0xlDkCtNJD5NOrSYnDHU3SCxOplP7ckl2MN1yJ+qc4t6aEqlh/zRyR3TmkjK3OSU+IHq
38HBTxVPCJSqExTo8vL+9sOczu5idzl3vqBdHIj00GrWlWzpjDIpDabupiHSRe+nsnHjcFTLRA61
qQzUDqu/bCCK7QtIDwTfRBpXkIadJN3sbn0VIebYdaS4jp48iGakw0llGfhfIME2dmqubIONDWk6
hHXN8uniFE5/CmkCzAM0Wqc8J/2o3/3H55WwDbuS/NPmv3SA8FJOZXtF8bz+sGjxVmlHoPHj/djp
gUzsnrJgohjymERmPpLnlytEA/Ir73XXoSBOnEMgsLVe4FlTm/muyp6XpY8tHT/xBPc5pEdw3yRk
L8Z59d43VLNRPLoHTO5q6MSxnd1TliBW6J5O/0tN3dBCRvHYhsfJhtE/gJYvyoAPfezee5smSE9L
7rBp9XXk7VXkYi3hA1ZSSmKpEk96ehZXGWbPzlZaV9Hc4CQhCUvkCUVAn2tSG3LzqAOnaCew3/Qc
1/mQTJXIGotjmyFhuYd0iMhVBrZvKQ8aCdNYv+oQhjDqB4FXn7WfY224kTeMsTjKUkuTzmrSrUHr
TcKtu0qRZH2rf25s1XWsvnDP2pVNlAHTtkWjYlQLJM+hXGXr0W6VkqY6jVRvrwa5+6ep/r7L/k/A
xlJd1wkeijLiH5xdBSV3Z3PH2/dA1yBqZT3+7refYU5O+jySEfomyFxsrz42a8CSLxrMWpwlOT0U
1sAzFYaIfVte5scUOoj7EUOR0ekQL08qCjV3mwlUdSEy3SPygiEeMzfvFBpHiQbS+1zPoJqXn2Eh
j/SOLHd+y3w65jB708eGFnYE3hvoPvthxOf34DCHQZ/yg7KSDmdtC1tJ0RiS1QHUvclOTtraI4bg
338d/K4xFcYSSHYqbB0IDDzDCOUxRtKpz8A6VfTgqZ7/Tgn3+KR+dvublIoO9R0mmjbseO4uTX7S
noUR52G8TL7IHCQnEGuGCtgARXhF+pCr4eXAdyVrIM8nkSC3NYDjtcl9Q316Ga9TnSb2WCKKpufA
9H1oKfKUguNBcvYcHNM0Ya8UNo/HwY5h9qY5rr0XnbYschNtsB+lIhQJchGLJh/SSHAJxfSY5XIK
baFG2kTctoS/AFta6H2aDZZvYKzA1h0l68/QM22peI+gg0hKJeCyoCBZkbD0UZlNPI2K/6BaPrVs
FkUNuLjXTRzXf6D6S5DjvIF6lTMA1AasEetkMUnsn2zaWLCOdPzJCpFUVrK/j5VyvnkhF8zM/Npz
kmn/R5zJi5KuCSV6IfJMnAgUTDYmrWOb/+STvzODbpg5WVaKMshvraQUysQHk6/p3eqXDziAgl8e
ubSapFkVAb/HVfwqrWcwCGnO6UbVKof+uRDcaFdxtvDPEwGhMXI4zw7N6ZLPDqUeFRWSRBb6jQgC
RsTAIbt5EIeypv2x+uZLejaqgQYqO2xhH7OO08lo4ZLGAHEonHgC+ms4iPNH/gdVIZap9CZvFFsk
hYufDSujdVxiswSeRRcYyv0qKWqPuX4ussskKG+dsizR/2GlipqlrIgqslR0hWlvrTXbbzBNf4br
eVJYAicbmSUrz7HvD0HdjA3tUNVKpdnoM2LH3pfkfR3ss+vIOgsvUooNGp7g1jpdj/uutKVRgW9K
Qp7Z+EeSGJ8kfMPgyvCFewRkgVPknUYkcqv3hfmiDND0kzv41LUjvwkM/vEWebMN9lwrRNXIwAT1
NjWr5SElhl2+oOXZWTqfaJ0tkbkZdAFzAdWS4GJsXKtHbGk8VzJ0itEXWOp+RziZZVDx1qr52ueU
54j0/XI8vTpJzdQCSOyYB6ahoYcw4HCmtG9y1sike8ImJywIdp1pZhhLB5rOZexZ9AR+QrsfzV3Q
qTAzTQwDHzAGlTcFJOktxc4Bgp0TbikNOOQygGwA5VcnmXgWz34YCwt6a8LJTxBKxlKM8rpM69qe
OSOj4ds7IfcFKCPE9FOR0a6A5Lj7/AXVVGpA/CIB3hizURSelufD8+/W7K14q1S5NxQ81GEcWDQs
KFT7i4GplRNIk2eDHBo/s/rSvzmEMiU5/H2aQ2yRxtWbaMv9UO4f4hdnsSVZ5QNI755CCrVzqjuT
IzyJo26VmzVE2pi9rM6UBqGonz/d4XfZJ7yyDMwYNai14zPEFuNsp2i5tuvDZyWQkZUA0gXyAPhL
6ipzETmg9Ll4NodaNUXxf0/O6pBd8s+99N3gUTuz0hzjW56P2Qbe+n3G3ec9eRUSQTJeEU0C2H5q
kVmgkKehQMkzUBWD9qUn0SM1aEbAv9Nmh1Axbs0ZAP9xRxaJwSqWYk21eah2CtruBMikAsuXCvvM
oXHrO5hKkbuqSqLX2jhvIjITr7RElBsmiLPcv2MTB6QE5U8VwQ4GMciJsZAkB/6tpluQjpoTxgF4
KDaQ4GPI5sMKPwq/+vZ1LHpQNeGV1R9um9QNUrgDJe9p05EHaBsl5w3gVvmfCrFIe3/vy83pnKGQ
pt1dCNybYRB5gzwA3vHA5RGypnerXhsaJqxhvspUGWPmXjVrU6du70mRvTxysxOEAVtQlEJSFuNG
1LV7n5ZcWKcDFoP96T343Uh09TerZzIKSNacEHrIcxuSj06N+WbFvSlw256WR/8Id/qVNEDQ7hsr
89xBCHZmLLMV3jVVn+HrTQUeRqC6XYg4yx/BSkBRPNKoqlhDyBNXpm1z7MCPc1ZdcbP/hZDjxcEN
JciME94uENavwaySLS69urAwUxI/u25+L482twyhofDnEG6pmh6Fo/Gmn697RUAMPdLplAX8Q7Nm
TCyPy9NA6QuGNz/e1ViuXMEhmvbss4L0zHbo2liQN2jqZUXT6aUV/mJUY2tiQP0fb7nvK4VsnOYh
nQBe8VJMIeVqZbmEV5uawZxuPRt+7gThr8Y5No4r9uidmQ0Jf53crb7MriqlQwLiR3bEqPTwOCIb
pZJZAgw44k7zboHdIn2kdXt8Cgs/QfJumrif65ezDmnkVFeiU9NEubw1MmBkfoytoMv3RepB2+Ll
vP9CHKv3hb4R2cIXO/tk8JhqU5tOSY4D6jF/+R8N16qKjl3jQ9YVuzwp+8QJ8URUjExcjvlzTmkG
HCzHuKDsXghsr0Y+qrxabS9Oc8QXV2f+8STHYWk8xJg362kHsg9wtJpce0mNRRs38Uxr7DCQQkYY
B1KdDKFnCUwb+Guz4L8LIfM4clfXCq9A7ajBtxjHVJNns67O405dH2VbfQh00p03397/G0NLiLfN
2vzwMGfU1PpBtOw9xvGWX1JKgVZ4ELw3ksFluT7X93dc2by1iY4CYFzGUgVUuUJYsxRAqDKug2sw
a9UyUDkPoOlH9o49o+OAEYaBotTEd3Rp56X1a+k2pfhx3SV08Gp15Mo+OY2EU3aSKRO3+3DdKYbR
vDSY6LVoF3BpgTe2Fq2pP9rvWrlsw8eMfWTaFHLT1meBiIf1CnyJZ1ey45ljAmVUEGmyGoc1Ljx4
YJcVZt0WPDH8IK+qVurrj0onsm+bQFihwAyoofrmWPjs9Q/qgZRqp9oggKv4atdGSdaJkKeImAZL
WUfKXEb0JeZ8p0UIf7QVLJ+10ozywL/PahPsf1o9OiQfoIVY4j1PXOS0LmCzAwNnJ3Lx5dAxEvRc
kxeE6f7s8XR9TvYCbWKyfj9JnTnl57kaDOYMUiXwkkOjL5n5dEeJBkHgKPxa2A3CgbruqM9cJzxQ
waksBubGidCNFw8bdvvOlUi2i/h0L1VFzxeNpjP10iIeCFnFYJIqCb0832dw+EaLExbvAXBE3wN7
mt4clkveGR6KrEOGk/mwYU5M6Cup5PlU9KjnOx7qqn09/UcLPqniQtNDpczPvMpkN8xgm8ABU+vl
T9cMrJICHQjuPSvHONqUUpp4F/2pheI2GDm9BHuVCQbePS7Crf5QyNz4WMBqGa1B6Tw+162KnAcT
AQk8D8pUXaVEnx+SAEKW07jI3ketHlFo0WLzMW6IV3ulxh9Yzn4sQklsGyRYugmRphDbuvUG6ks8
IKIig6llHOC2FOB8+B3D6BYbLGAO4Fgkw6+VeDGpE2lwA+DfBKSOHHqwqkqYinIB+jJTUkyLtXDp
KATMcbpEh0irPAlCKpv0w+ZyzOeOW3xN91jjwqj9MXPjkcN08CHfFSGF/OAGXkqcWgWgiO8fdEnD
a9pflsWDn18aPOROB6qQBTwrCI3V9bDNPM44LOnytLhK+WS7wnm5FIGKWK7A9k12DAvtemNG07b+
vmHo1uikEviPLukyb6OJOomw39R5DAAhGFWUIBUU36FBVwYifkHduFrsATiSJiYtcb5ri9wqFmcm
bgmuU8nmZDR8pj8HGpYl6eA+s19ytTSEFicK9IICHUv89iZAKc+peB+yMLc8Jo54Iq5mijYiF3Nt
RaRsc7/g4lqCSyAsx8ksvH+9WZyPWmCp9A+MmlnmL/xzKOIvjGekCUWfV/3Bh/egPAn8Apk0Lti/
xUhYWRH8nd4OT36Xm4VnGc+NaaEoY6XT5ZFkJJNlQ+/gc+eOqEOARzydseVNZzdRTFs/jkt1bfXC
huO5ZCuO1NG9MT3JOe0+aknXYIH763g8fZ0rnOSfeC4Toq/Sf/J2ZMCVloEA4ZPxq8QGbeAxO+Kq
s+y9cr5kfOMEdDCUzM1jVgBUiczWcy2jO9FEIQeKm5HnPwWvpeeAMtPHcKLO34vfm+NHexpiVw2O
MrcDTcpwAKlH+Por2St6QReZ+vKDv8lbp7wocFyoge9zFsz0vpIar0YBhiTU+g77nTB17TzJq+qs
T+/tQ1wG1rl9Ll/XyyUvSdXexR1JfK/wYO4I/P3QrZLz3GKbhbZw61u4GOgkabFRVrOVTvJFWOG6
CAq7tny0RSfR1X77Og0QjChcGMnKPVExmd1DggUwTE7pn2kWn204860w1vwiunAoMeo7s7kkFfkj
f6iJvz4z55dQ+XbT6LhczIiiZ4hjGLSZz7WUafEdAA+x0kJsYZlzulGU/jg/dNWSrEyOXQJWsryB
yolLFTBjIo7Y/PnEslx7qpdZbmxpuXj/WX1Tama/XzoDWaZo3qypDxEAqrrOmnKf37lhm2fv+Vm8
WwhZcfDEOb2U2nps3JAGzLjSTCtNJy+ZRPDUqhfx8gOMmel6geh0/MJMJq/4/rbthANhHygIslXx
mGTcTbwdFNrQK3CdjV7m/oc73ZC6UzTSIF5yo0vzr/A+t1A4YPMnzSSROisQy9290MEz5qu4tU5A
QoujqN4UIO/Uprs7Rvck+f4JLRHqN6NR+c/I2mFKZal9OXDLxe7HZQKk0XZr7/o9ND9DHDxefok0
9pyq2gapRbP80ND791C9NE52a7B4PWU4M0Qsea75aPz5VGOfsrMWFfb1oyyaATdcgywyjoKOIM+K
NVTh3mFYDAPpzHGZ6Sv6I21DVqSOzesZOvkUqhlOE2HWtBUoSuRtfuyi9yEilEeulDunCVlb3Xfu
8tbbJFZPBLcIRL2Da/g38efXnhhMJ/wlXmyhp/2wchQ3TcZZ4VSt8syvpwUvJhQdq4ISXYmaWBFP
Z3GaGhJogtZkav1fl7kr+fA/8jeV+ecyTCA65nZoyjKjqnsX93mPgnfk/BDOw9koAgFWPU0m3b4C
61jBB57cnJLK+kA+w1uqFeoJxUuMu5H7VL8KeEUZR+TU9J5LEKSj812OVW9khkJr4Le/i4vw+Ths
feyov8kca73CqvBdFiuhW7xoq1hNSBlQOZuW56HSy9qSNlDoqhaKZ8PmcluU/w8+UwLxYCy90+DN
xXlbLgU9W7HHPml+QZvecDgRs15tyIlHOZNJn9u64ye496ebXwlLuoYOPuifhXBBaAf3cfzA0jui
KzDJGBkOuXfQXu5T7taqXG3sG/6xgMd01PdI11ikMkfJXslHumvVZRvBUvUGb2TIxGlhlPbh+7bX
VblkFodz69flwx8wlCogxz3mZwfA1cYfNhkb3mlFVD5iL5VLnGsLvY5MpP6nsGia7n5/rJPfHc6B
MRAAH074ss6OA68Ki3KX+e0YovHmFC8WyJO9To0EHljRCnjPWBNx25+4raVMJynj8QIdWHvu6Xz9
SDecLQ7e+3IxKulVSdfDTqwFXyNtNgJWtJ0GVnNqan8/anZfisYplTfw3U0Vn56E47J1YF34wU36
p3Quq5KCkz1qrUGOwXqYq/YJkOUgIW1zQ+Q2TIJAkiy+pzYGgN+DrKOVY9sszUDZ++uK2XOp8S9X
zMjIudpqbbp7Gyny+PntTSh0cG1dYmx/VVBGTmrHu7CMz2UXVysRb9dsV/wdsc2PrABwS3xiVdiR
VYi6rbwUY1IVMLvGnAKRo88cgVanybgzfe52uJ59wxRl87Viotsj4C+ksgtydZaJgbdKN0AHFJrQ
QFcYdCl6gUYRjCM+hjjtBKCZhEOoy4HrT+Kjdr8FGzF6WAlFfSyJMwRauaAm+rrvBKCDyRA3pKCw
MDPsylgjFspUyKU6kzGjt/RqEsRA1HOxT+EVuMAuNTzSUt0hwcuDvpy7eo2PLssW0AWsJVQ7oLeu
i4aWNSQ7cGbEvb1w1/m3mxp+qgQTWrS2NK1e7d7eqakdVg32xwCZEFhBklZx/t9w31JRwriOS0PR
Eojd0WQS+c+UQkBeNKYihBDDdcglRT/9TI3wBurgdLB7UJogdwCPRSEuTWJTDCXvtRzV59RI+R6w
QA671DsIRTBadM5pbe3ZAJCbo/egbowkuH5W9Fm+oEo5CFBd1+qGfC8dRy7LcDNa/RxWPv7BW52u
QXNyXILoQr48tg594D2daxerKFRxavbSaNlspFR+9joF5ZNNN0IRPsS6to/TOhjcVktcXsmaIc/s
hNpjO6js0qZ3jsP4VhjV1hnlFgxf40mzO4Dyt7BG2LE+ka16p1tuk4xB0SQk3UOyk4CFshKM6QAC
jRccZikwTWUNK9H2EmFXX7CMeifcg7jBSRkdVGiBq1Bk8fdkRTlflsvry4FcngIm8J1hj+CnVBW0
937HmnQhKvKtQgjYQjg5YY3TzydUrGM8K6f7jJYibbU8j/pgMV7ZCXEaC2Uw2visKUx0LjqZ3wnS
FKnSrC4VP9CFvctqRmZT7M7TEC8IfE2Op9OS3WfoWDMi7c3Wq/ORt14icc3yRY7HaT+5w6oV572M
AcUpju1WY7uVRzRoIUWStG7Qiu0rFahKVFvObIFA7jPWcDYRjnNTPpaukqHo8poJ7tENG0wMauP0
M++7fO9gD1DfmtoTPtaF1Xijmzm3ymNBp2M/lt/H8PDgwJqFq1HFyr/4NTxnSS+ksEspSA2KUNCa
7PdD0OYLpEwvAHxGeENXDZuu9AVZyVBImOzMcybX84/2jr/b3lnxnjv4Vlup/GtrM6CwG8ZbulGX
Wl3bu9OxgPWQSbbc9rXyRGRaQJBxHKf2e91OH6XkkzuYrfVyY4EErDbLJVpR3A9kdjaS7V0PZoGo
SPtA6DuMczdkuQFuhPLm0XNCO+N2KUUzMwkqoniiPo+9ptIVdgcqjT8Z2fMwPhi4Q7gus+RbyJLS
EnVaXCcaItdnIsBtkkLCaVfmWjg2asDT185I7Ma5bat/NdLeGf2dFcV3bnJwsfVvqTkDGVWFy8OC
1wQI7O3CFNHPIR2dIxrAkcyxMItcrnx9lcRNAgz33ClPYomnf0RiX58tay5u57O/ooE1Cwalfmmc
Z2i/6ABAB/3/WzQBxV7Dj3NBulgEfUTmST2zvtJiISIp82mrjyfJdkoSqBSMmVX8thkAMSAsJ5wR
imS0crsdckhxmWJZtKMP3eESTPWVHxeSKRxlUv3RLxbQNuv1cahDZWDw1RZG/i/QYlgca79oSLYw
t41oAGERjuCm+DiUoaUtXdrfX2yo/MYq8RhO61osdCncuQ6LW9O36WfESYXSH3tCSCVr03LKUWC8
Ux7t1Rwa9xm6yxtTJ4guqsR0C1Ne5pDraNBouaswa1k7/XbA1EbtCvO1jsc37Nek6uPPmQQVK9+Y
Gmu19q+jdr6f81f2bk/FbC1rzMGj8OPwYjaW1XlCRT5ckVvhz9ly1IQVb6GjL7WWAZeZ4kcncsVn
KzzOy2wpzpN++0I04ZOHEZnHwKiWL5kvZ9ZQqbuNMcUVfSwGQxTDsaTXNtej/azTJQI7FEQ7CcLI
7/tvr1Q0MvLDT8LC4wYPGErSNDohVmGytCWgXRIDhvDLZb6Nmbk1f3SRONHuakQPa8RcDqlsXykT
6c3CB7sODXzbhQ9qnVCRsFuCLjUpQ+kYSNsnrB7tZklFkmri8q5ViBgU0YaBh9oMS4mBqt+3TuId
FPiay4of15E80K9oua8JiIo6FYAgAfZ5OoOOXsu6V6/PPTkywTRl5Rv3gA1sFHYdjDjjt5s7sMbN
bKRTFVdEh5AP9wdmYBlV+fgsSmv+mAiVc6D14SKm9wrIwroaw01MZ24fmxp52ywNJxIKgZ6N2Fsl
oG5QNAB8FgPX5xA9dkuam0VoxxNu4pruWiOAsw6Zt1Ajlh/qPGCVbUaHmoh13Ja0T7Jc78C4Dwdu
FPRohPOxLYBXXXeZwbxsDhJYWkdOg/9dCRqLlvxVLOVX4QURH8i9nr4dxWsGXUttzzLMBBX4AMZg
XXSErk2UL3qMb7lR0Iw2r31Ng8VeC83887c+G0wwTjuicP/K01HSJr2qH31GvfBxzkVEq8sxRH3k
d7dJE1+7hgkWUGqLXLJewujC1Y7SCgWJyPZW6QY4H3K2kk4TOEE0OmdoMNU3XIIBrvpZichbPubA
M+w4SEFOpVIOU8F3t3SR5WgI97eBbo21J7y8wZptvtr30bcrXYwy9K47aK4w3crNwTJWvsFC2P85
hkLC9zKy3o8YsZDiYyHeHJJ7EhvFNksN+GNQNBp6oA2ykP2cVAkGdXMi34NieVuoETGPBRxQFl0l
Z+hOTmx9yJIrqI6aIRFrXJtk1gQN1FdGvAtTJ0yWm0mnOh/NqwWixX6H9y+aSejg9voQQNTEHtte
L9yYItYjBX9qF7f9I+aik67Gvf9bGvGSaM/rFCuBBaO+9R4Z6Od0KPfvW48SFkASaNP/7A5VpE5F
BOyI7pVtJcqpBMJUUcqK+aXkGBVy+mBGkq6UOxC4TQfSWATxjh027whsz0AhAO2l3zL9EtSAP1hz
Ne4FXWNm0IT4k4ahaPeJI8cecDsqMc1G2rTw7waUq1xpqaPbYjioItb92BsNuQ2JNDoiab23LhIs
VUCrjZp2VnHHLcrlEXC5QGOCbGMXQD209yHMnyb3cUd0fAhT4L1USwDYT5flXhuVZHbqhw+w7pwU
xGXIznSxmHNKkQjUmIJvXXyqBsTGK1F7MGvjApDvyTBfN1RSTUdGUCIaScvsPpWYpJXoO6s6p50m
NKfn4E44/EZDeG5pKSXTMRmZsPcAQ5uRYYZvHgn7vc/mq42+6BLx/UE5cqeOcUuLBqafrgVLzbjv
LJTDdCej24cQxerXTlzhrOXXK31p0nz/ORuaMiA4DhLE0eEaoopuwFSdr8dtKWoKcxrFjh6qTZU3
yLYChsENFNmNca4ExgLTGscr9gLznRA9BpBQ/oTtr7AwkWINrpTqv3MRz3ScopdasSwaRss+sbIa
3fK1NI1loHF9CaIInima1pqIAdxY8va9jiN6V1CT3slVdTiLCNl2HEJoyc2YWcC5rMfZlEIWrlQX
Ij8dw/qyCRXqOzf10zrXJgFPqqBbImZAB9DbUmZpJ6cyTwar5UwRKmenEgsexnztnEy7OmW0raGt
xL7xfMjtaVh4Q7ekjGcFqHq9iyP+i0pup8smLUqscE1na3p+aWH7nI4IFrq9F1tPlFuRCmKEge3i
LECo+SC7RGO7mugOBpc34SfxgpwGOYtLfZA1L7aORR3mnifJh4X2gYZQ7hv2R9TYWDi8mrAkh0Ik
+pzE7ndXmXlhVCyTEvg3a9KRplOK+ESoH24Ou3BRqqiI4h7vvEh0JhYi23Pn4QcYV5zvOvRXkjuC
2A5ccoafKOEnRQcYv+Vs0osLcue5CicuIp7lYNvohlRDuQE6KfsHVMJp5hv9A6g0LHgRqvkJ/CCq
tV8fNWhx0WBx3bXqFo6TVaoBsk0odJ+WyAr9PVtM0/51IvpZpjtED0czb3pDtQ6uOnsW7aLSF0vs
zArPtYViCTWVWvYUTqYp5Eq6l+QsYLwbOYc2kYPGjcLC8GfvKBXO0xrQKVvgvbj5i6OoRXwOy03n
/SEaOXrMPPxwyISu1Fbe+UGBe9X/9a7Bu27pPqNryEPY8bVQyN6O4c+kyNKc7PU/n5imau5DT3N0
g8Q08B+QV6r5poi3iJrgzSHBe0UpwGXehzGqYpHTVdRlqLvxI9+F3G+DKN5W4zslFVmsvQ0rfVr5
TXdp7gZJ5QDJI+343HfJC4IFXemlJf9P/35VYXiv/yyXsJ/ibzVeOwkOQ68nmk3csP48HHsVvUqL
wKz9WYIMLmlXEp6+SH2vvTMEoO+860lQwToDMhWWV/IfLfgw6+3eNObW1Uyi1e82d7Bw8RHd2wa8
jVgG5PUHDkyo1Hs1DgzvtDsb6Q2I6T9ID3ELiHE61YFgzrt+QZFPgrxtLoE/H90aWPNnHL3yGvag
lZmccwxaRyHSPovVKlDx8YTwHEnbf8A35j9lMT0fklNNTzgwk/SOC4Ati57b7tBbHQTb1t3m3jZt
DopuPIjc+4Ig8xZDqmaOytcFYjKm6MVbaDUqULA9HB60fF1nq6TTEaQEiDJEaoDvVaRtjgnoKRTp
RgN2Qn4AozE8kmWZAXecYdCeD75rSNu8kPT9RCVahoCRaSBUyCfaWyN4TGcaswHYRUfxmeNCd+KF
SKsbny2tPU4D7KL8UTNyCIMapSFE45eq3r122C9DIMwQd3OBcVExIhLx/U5gFWwEcAhtJFDoe5K2
SZ96z1eLpEH4oD+VHS7tdpPifF2W4EFymkoCCLR4oPiZzb7hopsNV5+Oz1ysbOvVEqmaGx7ej5U7
txtSZa7Rn1BdOOCRU2d1o9Y7EJXnbtaCEzpl8qD+nGKq3PZ7sVxOtoGqch6ijNHlzrp8zhazZyEa
ZPGg6wlEOulGo99VDOJSatDVygHNGGktIPWNmFhRXsBUbXs81YTwoiRhAM26/CS2Az5aTnbtkJwZ
NYL24X9qwbdY+mrgIkymhHI6Go2NWU5yXZGqHuVNmzFkJ6Z3IaCwMnE9qSDoSEa5vuuuVzbYX8ic
oqVyZSufM4eLI63dDOIjVM9O7+29blWHgsIA33wiob8ebT2JFEGxT/hsE0lizlu/UbMYOu4o+rrH
lAvWVOXvKlXqRXgAZKyuxgi4rayYcOxEYBEXsrkpabkDnNi6ALVqjxG6oAFmW0KDDhzP9tmhNu/K
tgTcXtcQutncxAfD9A+5RDE0Sh355/EEnKtWrBTTG54rXGoNIx3EnMt0EBo+ZpCOvoqU6MFZVay/
QXHX+0OPNQFwbR/Wx7GtajMxVMpgI/Bc7CtxyKd4mSxkmu8qFGG9HeYFIhZoBKbcKnpEFGKH50Pd
Vf1b3Perx9M362t3/bLMW6tKhULG7ewWCSKZnxDcS0/zTN8a4dBbzmhfceYHRx6nmBUl0fKKUodJ
a5GTRUHl/fpHd1Ad1GRTaTPQ5p4MwLpL9gwKas6q0QdIoYa2woWXwqNiYtRqXDUWBnpYhW+b70ic
h3KGv/3hc78qM65H12Hab6Z2Tu21AZyogOsBfCUxREkp08vnATvai+NHCqKecaFhYA5ZAvtyiSOw
1u3FUMfBYlZvdOx17hjpgSUeczLpXx6t9xDT8C+/DKlmvsjC6BEzwA/F+dQf06mB/l0bwcWFPqSV
6NgutPa/wC2xeoB2qzKsxvWapIXAgbC0882CrII1xAzqRIfSadIa8bSpkoYhFAzaTs7RjXkDT/1b
mVww7tcyzMIWo10syN3fZNLRVSVCTtWPmjv1XOgvxBnQgbGo4DlLTnvg+6zAK3eR227DIwlyv96V
XeoyIbQKtK0SNISnYzlfbFQbudskwAwHqTxyOmFvn42nwZDazOq1SPCz1XcSm8T6sqBxdOrzpRiG
3kKeLSRhWddEjvA1iFCzm4cPHynKVE0YzWXXYT3JDvUQhjCXdQdnOxroVVXrriZb95RZf5kivVFq
ZO5UQ0FMxQR9MTNXBGV8ify5t5A/5LLY57dH+JXmqRAMiea/bJU2ZMRPmrxtIGwb9I20TTTbiE4O
82g3dMjzQBPIZYGo46fua6Og5qkY/S5+Sp8L39ToEDT6ht6AJMExcGJS2f32EDFdhYwIL+cAyQEl
MNvvSSKaWsJGbsRiUVj0WjXlJkKnaKLyNL6YGQKjgs9C8vG+wlS4Qu+O0uu9Y/n8DQ5xFlpe+ND5
mkvmpQig0aqnGPCOkg4preqaNIjnt0gLM4zJjjHELXgyv+XYKnY30B9ezP6HbDX8PVLzmuJCsSEu
1dpg2CjXu40BESQeGWUCF+BTQ4cPJNYgYoGTo7DvkQdF179ZvRqGKnXjCgZ8SAVU5WKHomFG1fkG
LlfM3hb2NQ8W9c4VNKYEto+E6dKiz69LftmALpgaHOZxOPlHgWaK9fNoTrez+fDrkuwgmojGqSmj
14ZD7U8y5C00RLnHc5g9yhCbPiGVk9HbE6rKWO//LSh7ybtvXz2AZ1TLB9/jBcFsioPt4Oga7+ue
T2QHN6T0tPralJt4xCnHR17E4UX77eeh1WmKSr7o1P0FBEUotp6Xdi5Qoh6Er8gi23t7P50NEL44
709TW2gGOFRs+U+Id6Q1TcLHvVBwJnsnE97eZLI3v+rwuGSdo1KsnOMVHzGnvsG5NmUHxp/3MtKs
9plnBmsxJnj4n2gJjFPY+7CCQgsYdKyLQ2H1C+3K0Zq2W/k3OCWsGWtxoaTQZqUsB/opX4HOFzk2
vlanA0PAm/NutunRLup3oYQDh4IQ8g9eVtFfVTxPjH0KcXsuQB3FoaIi+aGHADKjY3i2aDsH+12H
13ERwIepv9SVpvXujCCo1vR9wiF62T8i2KA8wU4nDEzREWtYvJ0bmX92ZS3Tf3fzjnTIznUax2qm
oKJIepzb0dgVMFqb8rere8mpMX/0Y0AO84e4mnJY91UrhAuRdJC+XMcSUIhnQAy8WcLXdQtQcyaV
2K658kOEMAnDeR/eJv080Wvla8d8NChR/L3fFNLHnHN4/RZsdegbZ/6gGlYxn4WSZ01fPKWnmkxD
CqWnT5f4pCNhyBkIqTMl+zpMv4LvLqC9A3u5zaj72CiNKb4Moy05l2iYM2hSuMHPQmPrDM2Ae+cn
mjPKu11HkLzRPVWX2WXEpB7ZKNnQvj87FKHQmAuPWuf6LLTe92Iztp8SfyQ0UqgaONRboUdkYjPW
QNGs2pxpPYroroZZDW+w8nkPgSwTcZeSenvzGV//csWwN6bV8AdOOlERYji9oa6chUYdmRKQwilD
aFM7fw4Jhu4FIpsmOz4SdxfnJl9p8OFopQ0xe451aTSM3uFaI0SN6vGVr9nUEb1cR/hZnOgBhQRV
sYwe9qTLJQnHcdiVzm1+sqYSXguzy4U5XLRcQpRK4pfSqnKR9i7mFIOcfsIA/NmUQdHVY/L1oWZZ
RvW0IV4eZ875d09RFb7Wc6nHduMzs3beK7HZMD80WhUd7iZUwq28EIbbn+PdU7tqumVInQ+UvP+u
Ryl69YHT5LbVvExgFtyYDf695gAG+cumsp8y1G0hxMLhQa5KTJS+Tnao1iJoXZRbv/Ip/LbOB256
wz8GETxnSlseV0nCmeMDj63Ua3LcdDjGaxObYpZildTjUE7HxjnqI+zMVeFJk69hJ9LULqqNeNTU
QI1hWs3oTi2NGQOPH1wSqmQWL8a4wTrRqg35eh64x4jUZDsC/TQ+3C782BEuQGw1Xjac88rO8mlW
SqtU7XYSB112hEl9FNEmC85a6J07jyb8yWnJDEMtFaZtduZSxEyb38EaL6WcB8xQ9zA7vyE9t5Fq
Q2ATYkMHPU5P5SnAKT2okb8LXtgVEmIIlwslqqdpE9bmsB49noWTO8DQtsBSb/mXuzq4q6x0z/Y9
+cG68obDwML/loOuzt2c29BmW5yYIqnn77o5YsLH4S33bfNlJi0Kzm2VgqkFClGPTOfwkiApxNM0
KzbY9J3tbSBv7YQwy0M5LYTO7DgkxIsQ0sOziOojXua5hGtLSS4R7sHdn2OQEA/bWrhaMPyMsk8A
d9cgnHbhGhOEhPDKdUkZyFWJpPnaJgfJoHTGvb4fXTQRiQQctOHSPngXp78M5MHB0IzKU/uHhiQ9
6T180resvgBUXYyrhC2RfJRAm/Z6M6ZnauZewL03DVjMr4UTGclFhsE+dbNV6WVv3jK2uBE4Nsye
6QvoTRlo/Wq/DULYdSK1c+DlKdiRPryjNbmWBep22HM9ZFDkE4kscUAKQc0obSdi/22EAfcEsRM7
mQd8s0yTStvAJu6qznuslUajkDQ35EPXHkULLisZ6J2i4T28zv/EwOq/JRh6IfITyw+C7hC/fr4w
oqBu7eDQyac7L2a1Op2hHVyDhboFBRzvjYvygPfC863SD2nocp3laXgBKrE7zi5pjJPiEaMufp3P
ZvtZ+mIHVPJdfczfkXJY4G6GNJxPqbwWg07pXSxf2QDNDs2j7yslgDsjN2fnYSlsR9NJAQRXicwZ
bGcEej0xD1vwtPiR6P/EroxkR0/Le0mt8i2qOLD9Rf5PcgtSp8b6at361tby8/gXf45L5qQCG2D7
s0i2qaqP2GpXUrl6wP2wxyjfEExWqJDvBANNi/sZM+1+kjR3noayymfyQ/gPKfC/wVSw+kIh+Y4F
rWeBHkiddIRn5H4Wgb2/4nx0Zd62cRAgya6++LvXUFtlKUnacHgrUWOQxDU2Dl7TqHXFh1+8/+Hd
zixCIR4SdGHcGy/z8ZTIc3BM3dPUZ0yl88NisqTCatvPVABpDqrQ+/R6Cb2NwlPBSaRj7YuCeWyK
Gngfx4eQFlkH27qVgXBshe7bTx+dfE4c46cn+pbPJ7Z6zTZEnw3CK2Skd1I4B8h1Mcaj1i9iSNpe
/kTpLvWoOXB+kwgivdkw0Pq4YdfkDIXtpKKSH5yodPhCw1o9TwKbcg1aY3LgfmmBqK8JBCWd5dd6
orYpc0xlUb48AeR12rlN0mMidG54p1BbGM+CG1KKyYLe/XTW1ChqpYFNeWl1hVhsQvNLSuermEEm
8TVBOMvqOfPhgGGrk6gl7hsKBk9uphORp0kJaBpCSXpyNl3c1B4YA2t62CRpSdOvS0PvWdfTJojb
+7F9kiy2/fzq+pRKArPb4xVmP0MJZSuQFyhhcx4UVzrD9tq2E5YghsnnSN0kEqstitxJiE6Iib1g
pKE+ZD7bLlS7TC13l/BSmUzsTd3Et0YdQuxgGQszh+02YBu5bF299UgUFolC1F67ZI8KRFyKMF+d
OffQF+hOTtndkXnJhUA6bU3QZakwGp6tJ6gGu77beN7N0/TegzM94wj/5wWs52Q8/bXCvUaYIg7+
Aa8Uf6ZwOZ4U/2cnFRJH4o19UJP1dr0fv0nDQpgTWDdj9gC1c9nEeD0b9gvzwpS3+onE+2mW04IC
D9YqSKcR8mzfbauMk2eTk/e3gxCFV2mCdocn9a5hB6+c5t7xNvnyEXPhd1QNGEYll9EiQ5F7Eoud
PtcrcILXumArI9GzvTp0novTxQBLA1XfUVhPiMNhUNEBGdpb3s/jlDGzOTM4b+D/vcjEwlimg/GO
qPsJEZqonys+2eTl/Ov466PHKiTdaiHQyx0KdcHNrIErlHwyh0M11inb10GatQtzrrOisqyaIHnd
OY0etXwKtEsJX0b+dWjelfUqI2ZNvnEyjuvru4BMoUhXC8uOS+T25tdAnFfmXeacABAUt3Zn1bFC
5avqD8OPeT5TiNIb+5oLV8D7rNijlsQ2hwWkYls+Ce0nn3Rn+uHhQWEd0LaVpgGRWM/LJ6o3IkaI
JeoVnZOP+0ZxeLpCkedyFIw7UJo0NUExTWWc4N8yUz378BhdsAG7OJe58ZfQJE+FSMfymuLsMZng
+uMnGcb91y9JsqUuECoH//34330j+MLe3li0bKhFeLCrAKfMf2td1YOS3ocS4S1R9cD36cT/juh2
YiqUX6EFY/XU8ZkQ0BnN0cGiuRum1u6DT7juNYz3GoG/beWuNQyh+Dt2J6oOVEVcZL7GYWTMqwfh
5JO5UVdMrJmr34AJQai0COSn6csO7CfpI+ldxh/dVdgeDR+GgxAB0AdnYdADjVYPsnx99/+KXVsI
Ge1TQWdVdNc+Co8ndOTRAsdxM5p9AJLi8SLJ/y+DKi5a0qatRyz6cu9j/wjokz0k6whdLLiS+vAs
X/r/gk9ZRF70cGWWV0T+l2pGx9JP0bSVsZM1JzrKIYqPBRWr+HZYxWB/mcR85M1vPNq3P8Ygyiuk
QvqyK2kcEMB05MoA3hW/PolnRVCZAf2aTD2tnHd4Bop3Gw4I3DVhtmymz8IcvLC0fMk5Z4nnwgUh
eyXYFFL3xbjiG0t1MoYqfbP/t6YU5/RzXldADNyXS2aMaOtL8GZzOj7JbfwMt7Pwa/8Q0xepJ6AT
5F8A70iK2NlakZ4leHCaWn+vI3AykUY8o9jANqkP0/D/6L4E+D1ql0Sj33FZCdjloxsoNdEc3TbJ
fItyhgSYU2z3e7lP8QpVDSImZp9YJ+v9Ty7YBkKhVrCjwNfdqK/RLIHF2rxDSLDTQt8jBtDw2nDJ
NHQ7x+C3fqjbSh+07JrHqbHYJuQUtUolnvni/5rvtWYBN3J+epOET+HHPk6ZnLobRTxKo9EIltpg
Reo1hUwmStHwD1/e1RkKgecnzDNXGfkvqED91DRrs2RXRRG5GdYPUQDciJqTEU4I4V1+XHP2c1tZ
M08J9BC8DqJh50AKPqZhfsaF1AuAj1I0hnyl2optpSOL5EhLgVHE8gmmotH/7ntBHeQ1FR7qpgRp
0PmGj7Qo38D2BFatdFLerWtku8tCV8zr2RHhstHV8wmrCCnCQ+14lcWMVVVF/cXtw0J39KEdT3aq
OtHmaNg9H+Go+pKl0vvTMfsE7dD6/NWsAoKeCkZ5ppqI0hnHZ4PTw+4elA/YthaEiFSNCyCWzNYg
hcL4fKk0vSSCKQCHU3igJc6jF9oH2mT6tPFRE05Q+Hn4bd8kcD1PohHYHG8fjOpYy/DHiKy1Oe+3
UZY319tvimpo4r7DgArSpMWY2R556rU3hCfkOT1Jxsi3eEyQUR1CtOGEgTjpfx+X33CKtkOoSYln
65oTpvz0Z4qiHpb32xpq51ZLX5kzRmjqCfCjnGgAxBcRZNZR6k9gTvP6SQCkLEu6ehWDDmkOg6k/
7bmsaZbTriDWKeZLubyNAx2HdT5R7SiBYwELIOxQZXwV1i1bOVzhMYzF+JrFOSslVwgxh4jmB6OA
/Sve/SX4haE6hcSqV76NjaH9zldwfom/oS/FMwY2vl7eYnM09x7NCqCMrX2W2n8Il/MNWaVYjq7k
DSE6APhI+3VQMsltvfgTCr9x76Yzf7YL0y6q7PT8QIYg/+n9yyeJ/bM+jrNOtF0VYunxn4sp6C1r
AhaqOTpXjoxe9TBhlG7Bq74IuIyV0AJVvY3+2eS03sMTMyyrPN4VCIlP1HSgGXbvxllxdXLB1cjc
EKsRDIZ0hTyAkEO533BfEf80RLCn8oZHqQ0kpwpncpZDMJbmH9F/fQqOgimR04deK7RUWfdnwUc7
WRQaE2c7j3bx+IE2bXyL2MpHt7qum1EHpetkF6SGZ3oqTcfKk/wQvc63lY35/Q/ue+ZtGAzD6FFG
aZExQyxjvxJgUEu+cHdtRnGT9RQmS9oYZXZARK9KAzN4TClY1jU2ddyXRm5FPAn+nnOAK+5XofYq
j2O3q3RO2v777TToymK+AvkmjV4b83coDs20aPOBs3O7HFeVNHmf0ObwYrKzorQZMpLrp4IAt7Kd
qWJpM48OHmfAdXIt9313tzLOFBEfW2qu3b/4zo1gz6ZHwAZENNjjc7jbe9v8MI8O0Z01xFman5Af
PFrTtCXKo0nNvObC4cgnEgTzvxdrj6KHodNLF486eq3MDnjigD/bwQS/X/eGCu+lo2PksJPuReMO
jfIld2+1ias4n112x9+zOQV5Oo11QgxyeMF04nRpidi/s8993wSEhX0FN/AGO4OEJrDICBIZZpg8
YxnFA8JcRXr/H4Xag0XgyT6nlcuWilbyDmHHkMwo4BBYe0qvMBDAu+E3vSGIeD8oCvzKYDd/jBWf
jvBWDqpT0mv57JfxHyhk1IaZBi5VBE43MFB5Uxk+H6OUsB3Jq52DqKDfKkZOnsg6jV4UuawKoWuX
c5Uj8T292dxzTt4tg5qhPM0FhgxYOliZKXNMoae9ABBPPHsHgO3IDUrZA7fO47hgc5X6R1aPtnZX
YhYc/R7/UUjZK1b6yAYAKpuVGIyCgsqiJ5kblnWAhGGh4x/ny3JR2bTY2F/nlvMIwdyROvglekFW
axr67ZgPULfZhq8r61mqbBS9mFDcQ4hpHGcOMJd0SHvJsDdsrpCmULJYZLeV4iYTRJHwf9EXJQEf
wW7ho521SlJ81+tkVPPEONzugkPGi7FZjiqAAA7088lDvTHv2xRAS7syIsugW+QnJSMrkO3sO6Xt
1+H3DLCmVyY/ytaR8s3o4KQZQsytTm/kY2B0RRj7NQW/X2pf121WlSnz/kYm46Ppmc/S8hFc+jWf
Rhranmi9C7x+pMZmQcvxjFfmwKQtaKu0ejtnGS70GvFjUX93lIsdxVWnIdkeLN3ONrrFmGBLzTcN
/Um7wYLjjmyLL+FuNjx6GBVFklsVYVSqyYZpD5kWUYpVMUeh2FXviLPn7rbf5RQBFxfOvyTN4l4B
milGagWdkOGCIukJeLD56ao+ahqOPmK7kY33uFYuZBWQ0hM5+wMkWJAgnztBTO+tB8Tt7qoMihLC
LQnecyx/Z6JxLQFwNSwHF03Du7uJPoHapjs6kr97UXuxW3PNx0gRmyG0o2Kyll9K0AUIhM4OFirk
6IsHhqzkB/6WJcbiw7CpzyLfIevmLu0UktaE2bG+pqo6hmnFD0fUKOlOOYq4lLB2cCqb9hj88UKA
4hG/Ezw1FtcSkz7fSNSX7zUkCOrWFpJXwkPchTp8/jAWfsZC3U1AjbvH5zOnOXCsyDnW6MyYXoR6
yYBwVL2Dr1LcnMIrEo79rJyiqLJ846X8IksMxXl9HBPpwe6qwY40zFI+v53cVVBsvyoB/PSX0uZQ
XSKYxb7uITRVllJFPE6lAwwhNTzV8pv0Dn6C0fkIzDp13Zx56LUTpTJLf7eBAyZfuF/YCH8VRU5E
zbTwoSrJRMxBJFNcpE525qWJA4JELdh5iuOsbB4BElnAc5VWXPJywzzW980duf5UxE0AKUEJ5JVH
uzI5oz6o/bOvoMchXwctnjSI+Xe0rENq3f/6iHTFG6wuiQ8e2iW+OShHBDBqwZghVMSWLi44Nya5
rv3L3qQ4gDMuUND7nlkz0+qstnpzsD4ogUYTl2RO6M59Fbc65WTgPd9GsN8jfam+8/bKKcugq424
oTNcjxP3ufiEVqwkwyXZexldjBxg8E93ajtxPHlBDWSnSnng+qaeudMhY2ImoVqw2opqL9Gi3ZER
Lx7iGLycUIcfZ9lLoRxBjcNRf7LoBfBN5EMmSg52KcogIfCjgGlOk3M5Bmdy4lMgdq7qFpR1BGgs
Y5SXY9qhKVHzvEe2l8fU5fU1Pnat0+3uDzILUGWUPxD+g9TYqKMeVkNCj6SejTLDkWPpRLyn4iuc
kUDKqfVZbeOLxPypqTL3u/28QULiuuVthFvSxwWJGZLBqniTHriM0uTOAl6Gubg7f4m2v2o/BTVm
tloe5U4O1dPioAdBEnL47qxGr3FNB8huqBTeGi/rXEsE4kBw+zj7PGV4rGaeISr+tyeLE9VhAwlQ
z75SQsMldN17gpK2tXlHo8rIx6ue007a3jEO511jV/jDG8BSeSCUVdQ/0z08x9rFKmxtnYsZTetf
ocoi3vzQOLnKLYkWDQJ/l1AGTSF0QLrNTsIkokFRWIxeDAKuisXQdyejEo8Ynd7euwgp6mdGCTRR
ac/OCr3MC6GcisHGfdkSGhfFlyRsRGzk9lM+qM1rnmtX9wqxTFPa4OvleFodGTkaKKQ+wrf61N8z
OAT62Tbo60SBdduSO9fnpgYsk6HMboA15HFhJLUBUZKRupU7RSOY3WdIDawcZSvLzj++MtB2dRcZ
sYZ+TM8YrbHyrJfIFG06mJ911Ib2NzSchUIgTcbFIocQ9+vgsD+ZoK0Afp14/7ik974ZJOQqrSOQ
9N50rE76jfCQrz35/dPIlpYNtLekd7IL0XQxuykLbpxqvBkbVjbV2ExHGzjWuKZpqrBVB8m6y+IJ
nRHLnSuFbUwKv+rJBLrYup5BUbh/p3cO6grbcp4uB3eOvJ1/FfLzqWrw4bJzu+6esLBCC8tw+ABa
IOrmPKyKr9Ku4RHyFjoJdeEQcR0+9LrGd0JT2JNn8cZhi1zqkzeIw3oaQAzlnOCDy5ejZ2CDfMax
TXoH56lEg8iyNMb5a/LyZx0QmbcCvRr9fuAFD99RQS3pjlGiV7g+8iZ0yPISQYdFJnqph9FqBeKq
4++rr1hJ+9hTyN9DPo9DkBZkFZnQtF013uOSfShp3lHdt6Wl31agPhEIdNbvpsVnRcT0HGvyM13c
jdUnu8uNF+tNUUQK1hlIdnVWl3d6LnxyBrodlcgLy8svaefEmUU/fZGt2LHb9awIhxR2r2ZsFIHr
4Wi6o/26VAqRBL9vlgebbhaLRL/T7mMI5EgU1rFFVEb2B8p+7pFURfu0tyBWPXXBcea97E+TiPSA
GNcTA3zlsY6gsduLNvc0GRaj0LjUwltMK+nOiXyYop51+0RYE6b4i4QPt+BMuD235pY7B9GpPJmY
LJZQik6hTi/Bg8NWOgqcuXaDWPwqL8DMuCJctOn6T1gGLVbd4jXvfmJQQsd9XF18+vArTFP2Z24g
z1W4V6lCE9UCN8XC/x73yzHHNjuKWKLwEjuFNpyH1R4WnW5I9RsuD4qx2y1y9am+KY8br7dLY/2f
1CTPBU5JPIvd9aB11+KCvcbnC0Gbs03zGYShK7En0MeNbX1sfb8xy6AzSzv8Khj5chBfEB3xIokb
Wujl5e9j+jghcK3/WPtfRd//E5CpwPzWtjHyOjC6LNaS6Ww19M3L5RDRsCOnT8q7dCm8AuNNhveZ
x3KcV3TrjwvSCh6KO8b3HCimU9HhbR3NeUwOohh4YbW7Ml5/kcLi9I+aOywmDPjlePDGx8uQeN3G
RG5/dlgpSDXc2vpxZKRWuelrq/nicQOR5ESbn8mxVJZyQ39UkKaHgs9cJMmkFzlkevSAqeaaK+YQ
VCM9LheRi5jaYaU9kl5vif7thnsX8m5YhsvCfT2/sT+QFcstaz79XxB1wfCicALubw6eHT9AcMJf
bfrF0OJp/y7OBKvkFP23bvpaRf3bLwVNAL26tnSIOZk1tpbPeZdwOg6SP8I5xJIuyv9Gw+oBSDgl
b5K5h519Qw3mO3BRHVbLvdFwSin7DFJDcK16CxYpq94RBS49ePhWvz6BAs9OTKzTmNa+m+3iqsRQ
zPxbXDjBPMWbobdHDF5A5cAPS8mFyuOyhnm/k7foxhjKfXiJBq6tMnBJwq0+qIHxML9k56y3UVxO
KFjZ45tN16l23yrsCuVS8HN5HaM2jHLIf0RsIZA+Ew2W4sHS12OTCvSRgq0nqdlgzUrFlKOs3LZg
SeWDQjfIGHse7DgxBu/1pgW/GH9CpwIOMdAz+fHtYScw0MHU/ZBlSvOz4w5gHb+wxwuuqDsYHISA
OO8ID0VvlaOZftxkckEOlWttzWEnUSboo2nFnTyBMs+ZxDPIDGHuszWLXUJxYBEI8SdtfVTXQUzs
ItXfZT7p6B+cLT0z5uaJRUmHi23JfV8fGjpbp/RD7aMPJPRUhielkGJQCT62LFhnEx6lWcygiSGm
EWyZcMorYefMtDWi8kvFJUiss9MWLC/qPpRiN/5h9vdfSG9FhgWprqMxDNd+X0v22psOLwfkeSYP
iOWetejVlbYgpDvT9XQ879dGbKyg9GbuQU9zashsnotXnf0aaEwiFeXiKFvJ0yLduGs7W6fIf4uP
gRvR5dRAvBwojAOKINM8FMSUNF4kAhZu5CjxZYuyr9SxLnHKV5vMW5QPqNZZ4ldKIbSp00x0M60m
ppaxpAu+T72suXto2GosC6cNJ7MzEDIUPGAcSaVWisjBt5XXd4DjKtfAL76l9JLZceOTuwUhY8ba
xv/xvebDFnRrN8MEYJreFGzz/hSh93D2P0Gexb2EQN12s3xIftHo06ZU9HJrxn5wtHj8I7+zrx1g
minvV6E4pWCSPYO11FM7PBf0aXKmBfsbJ6+VNOXn1uqvTtMqKRCc9EuAlOXt41OkJ+MOiQnt+QW0
dkUACDV5vdAuwUEkG5daeJkbBrPDu3cRVNkUdk0+hhNRK3nbmx+47JYFDwdyRKeYOqqxTfQGQhGm
b0UV7gX6eaLFMe/j/G0puOZVc9PkfONli65XSQCFm3dXo36or6Qb/qUVFXbg9gGM9ZvWH2JsB1ya
kWfBS3BAbhmjvBlbb6IjlMvtY0hi6eJy5KJ9PLymcgeu7UTw38oy2J5ID8c38AgUIGSy1bweZ+XL
yM8AGoRGpJl42szsM2G2IcULMNraZsYHpow5pxE0hwxKZ4m4J9FatkFfkZVOWNqq0xfS0dXfOj3u
X27d07jVx/L/gjv9TarvXza6+MpjCJY51iJ/uDpxgHwE+rCnLZOUyzQxjAmCU3he5yICgAOuc5N5
hezvQd5Wubc9O9BMiHpN2r7plpi89kL18Ct5jLz0lUngYLkfNCHw7RJdU3yN71ndcLog8LOgvfM+
vGYeUy67CWCLuxbM/4ekc5jtdiHAytD0SUZbkUweu9veSy4oCngLVN+vqK9zVgIBftqQqicwf3lb
1ZHoc33P33Ct/FRVotdC630lrSPo/eLhv8VyW3TdbS3zz61cKSXXu+nFXfydSqTMe1SPhJTd4JKi
Yxuu7IjTXGtoRTgkbWqcyKRhlZG9Nwc7/zanApnQwIdvbzRzhvszl+62qYnN5R4qRMbJErZlW36d
PtWrTx+AUBWZFj9UjznksqwMbtohrPOdWY4d8BePIVGTRpiBKEgSGIt95ht+8B6+ATvXhPTPjF6B
M8qAiSeJkX3t2MsmhcZ1PpXt97WMYuCT06hPcQss7eL6jSMI9vevuLvF94gaZSV7UzGSqmx5c3Uf
1fEXxyXxPnnUa9acVdLUhrl/3wfS5mBZSaEVCp5CyZqd+W+H8noQvQKwOMeeh6tL5gjAYK4i9Gd2
sGFMor6NBYPcdoIhuAia9Fb6Fr5to6smePBuXwuD8Wz1WKBCvdBQxRiPyWAJTnbWnMTE6TwE5yOF
rLfoVE4BSRbJ9oZZPKSQ+WiRG+g2lWAeRv7fRkTmL9l29G6RBQ5xirznOG75pylBta4m7so3jda4
Q0t45Da38vDnlqh07A1s29tTx/G5muUQR4RHPaIbCiOBJ4DK6Syq2xAMISw9DnvRBuHxKP4gQ6rH
O44oCKriB2jVs643/gZMePq8ezXl1azcAzJuF+qJD/mTAxHmDZsmSRzmqVUB2j723DN5aCbC3n3C
0ISIZYDKg4LGxQmbOrPpND/PXIGyTH8YgfsE5T4Lokt3borM6PxZJeW2Mzl44zrB5TYWq23H5ygO
EhOhaimiz0Lyyb6Zz/ddamikCYcH50ToogBAjAQcmEB344H6n9d6mo3N7xwCns2P1QJOesdzWxva
6ll0zYswcYlgiz09ltee+4u0l+1z/ERbxNYspMyHNR7FIW3QfeVwR6B0QgrcsJvqZHb7VTWIrKyC
Jza9poFtOHzR/sduBCp1SVHd3TaK2Rd9ggwX919koFXns0Y2JH0JIMYKyissew+5jdc3cygH1p3N
pkyxzBAOr2wxS/kpcAWaPDbs0OvbMK4K0U6DGo6ic+Ge1Z5TZPOfUSRTnVyIjdUi/uRqZylEjudE
lSK5ifGr32JLQIO3/CsaDm8UTT2U0WW7uae/O+FjupaoQ0jMWmx3jd6pYypdv6dkJUUpKPXtmgT7
uvXJffNLdb+mDnwrMLaFkcSlXIONtXu/T2Q0oAUsSDdHp1ci0xAhx7LV5KiEcAld7muu9QyyQid8
oUP13VhaXhLS37eO6MpyMRG0vfCkfwBc/g/iUOr+HsH90IHFpJs52qft+bERLqukamGQ4x4nDDK0
x5ikUKLfDQl6Je8In7NT9/dCe/Ehyrj/2hb3rle0o0g+rXhx9YQyiNseDArLVYGZK12rhz6n1Ocy
MDolS65hwSIgeJqneE66i3NfhqJo8HDuKlRLFs6SWzbbIQgG8toAaHmLrEQAg02oQGX4PoJ0dNEI
aiTWQ+UmglKHVjQiIGGiuMYfEsqueRulElfmxe1AVCNM3uOd3DBesRUMFcY3pkOLVffwvUYhDOar
GdNehHoR+0/5AOJScsdaE9o45y4+v/EVKY59JxNi/F3sgDxA7JkCoCwDaWogKEGzxSJEa8uyUmT1
iYK3dwzRam636JM2RvIZIRHzPQaZ9rSmHJbENr4Jewbd2XTaqphw4zBUvazNenAMxswu5uwp7tJk
XeDjUgGk7YQh/QQC9FsexH9Qbq6exSxf0Nv1Hx5zntQ/rMIzmeQLAW206MSHCAGV3jDJcQL29954
0DMUIEMZFuqtLr2EH4ZeJAM2nTE0j0YCs9TUTKg2Nt4MOI1JTH6c6+4aok7SxpV86U7+nUz83k8n
SpsaRsZ9dH+He+ocUJxbtOLTvY2yhLEe5XIiZfZ3Kmep8JoF6QbJSlVZyYmQTMFbGAaZmStTmtRT
81GG8s6fcKD1qxsaN8d90cYf31Q3J8f5BDiNuxfOjHN1zzX40LSC6CtgoLSjnr8XqUxS8g885rfl
ns9IWVAZx+9QXbXQc8TxKFTXBdMrXVEnVCdudbOBCyZsfI7lcnUzFSI94Zn4peGa1rRWQUSRR31R
vq8nOIZzO9dWPYZ6kfTOrVj892+8AfquBG042eQBvTTfuh0o4sL/Gq4wy3qN1/KUmbBI4voAdFjr
yPhoXzrDoIW9DcFBcp2H2c0GHs2ExdFzZXenhdPewZTot6aQGBYFQ6TAuem1DyvtwtsJfYiDvDzb
39F08/vQzh53pRsYuDVIQRWodaEmJnQQSm58nJyDWClZqhCN1iqOp7KsOiLENXLI6fRRmG9gg9d3
iiCZ4rpf8mk5nhGHStr2oY6MC6yGSRtZr06Tp9k8vxyvDZ3YDuH4LSTE1QhqIvj0dHXQcG0m79Py
TsUYnSj0N+8BwClgBadwrwHHKSLMCdsXegmR+MCt9lM9raJMeM9VeQPiMXLEkMkKLc6wojQF84IJ
m3t1SII+Ln3G3Xn0FLtZgVYA4laeT0dnj9CuxIDfGhfgazS3SgtaumryAC/Mr1bKSIgQmdQ84jb3
xsarnBpzqN/IeYxwcyG+ACimEFu/Dk+luKRJpYSDqYNA/ZlHYvns3qj/F9NgrvM7gTWhOU4pHSfO
ruedOutXl4B7mU1Ts7lYvOBxorSKdeffSdT7Se8ImEH4+bVP4EvSZzRgcxj320/z8P6QM3KvBqli
eJ/W6D7rHZ+KceUuHnyDs0tBN7ZY67TwN7UdVUkNUubUL46+PoSZWBXG9FltkNwBVpHIS1fo7CER
+k9Micijc1jpa+qb6Q0hgigdvJcLAQzPVi6WqUxRtWTWrK7vaoht8UnFwgHehEuyspNRJKNO8J3J
xZ5pcgKntCsHDYSrWC8lT8gnO2wkn7u0bG57UW2qLLA4oY3QqrXaRBquYLh6XZUaqmOsxiFcU6D9
aeQ3E8RR+vN5vxi0LkdtOZTdSObUkrvWywuaa0QWywbT26pZCG/orqC97NKPCG35gma0k3qdkRa3
wz72zf2SuLdMmx9lboxReMDoixF89Cei1bROpolSG3vdpnnEnci/ichYlBITtlUozicxoqzsIH/c
Q0Tc2NYILvV4bQWE0yIlWYYPxRZPhC2/plnz7kya6NdHTFSHmsOavjtv+dN9FLQTgJmC799Xbej1
ahpb2xcLyUCZKBXNWaheeMUvWH8ZfXq+UueSGoNV41xugn0SEUnC6yhPyD1OfkG5wyMwNVct8/sw
wL3XWvlBOCS8wyTBQtoboU/w6kS65J9GIdo04X674h8aeAdqWrOPOz6WoMNuA9PSfC28QHMEDQFT
AiG7DJ6Cg/z27jbXRcNsqJULVPmP82JxLjqo0ipJxZiCMhGmCCn4Utd9f8Hnvip4n8TtjbPtaHxe
0ST+J75c5Mtj/peAFwtYhrDIJFMu4aW79MBHHbUrF6qILQmnFEDDYJXcM1uO1q6H20jLelyLt9zq
7cNEP1TagKHN8vH5KC+YwzenStIfrDka2dKj+8eEkMDlT3xwncp0m4aMWA1Fw5NFGSh71Nio/GFy
As70uYIwbDM+2fWxoZx4npsu12f69RJYsS7E8S+1LxMwVVSbQEB/tMXzMsEIxbm70R4P36XWHhcU
YUwCYmXQVfGNBzjrulYjaeQL1+paWe3UqU/+f8ReKXgv1ArIaDJIEQM+gA+YP0wplWeGmfEM5loU
Am7D3Kwm7biDArPyw8Zen02e/4WgWNYGmFsyVX+dVP2bHhcFVCrMO78o+u9NnBX+MzbdQ2/Wdby7
7Z3N4V1wT+qNj7SIMZ4yn2g49rtxldDbBnGD50Iz2NduDb7AxIdC+ATc+ACjKPpXzJW4cgAwKunT
QsWNsLH7A5ojOV9JAUxKtMqOfgNNOaCuKy8iBfZrXpwvecD1fP+oga/vgS8rk3Kl38j/eDgKd+nG
kgrYr8wtnqDm+esw4+QwQgdALswfR1gFCYRo2Mt7N5AGYYS6GkYtarOVGFda8SjLWX8ZGbLy8pBO
9WDOFdhiQGfBzOf/J0ZjRnjeiuuJbUvOhyTKKTAL2Siqby5gmqrXf3g655QXCM3aaW3OxbhIjZJ6
XNz4UTvHBJWCwQr+ZdiZio8x1oK29gjOcIEsTGHo5zYcdRxERz2pKrfExz1e9+kjZznzDCBm39aL
8Oc0RXhYWoa6uxwekJYMjTd5FE0Yum/cX8r91zozLZltTacXmgbzTDgXq7K98683WbbnyXRXCQU6
f1RScizycUp+W6IlOVGr984wMrqYI72nFKaxlsZYKA8Z8po4/ZA2yARFpYk8BgNr/9Opi7MllP+H
5aVXyFLsxtz7EGqLA/6t/LFWgnE+O14FGnWKQzSe6Fca40wNtqqI0FJ7+lr0FtsuATeqQWv8/W0F
tUbvoRaB4bBVd6TGeMWfFhYh7b+Q1XItbUy9qXOpRKBhvm1BcETuXcbFuEPDCRtoJX0lO2sfdYOL
J+9Z+BsrlCpr8FsLKDDQSRd5Sa4/pYJTyIu5katSzwiSEkuN6Jbx42iM2PReUT0/KWKZkvjWJEzN
4taWRBQKw8NE5AwUg/B6fXM73IGw7KcYb1x1TvHYUGR3hLO9Bm/NWlWqF10C1GfLpINMKMAcKIJY
WF006ETURUZh+T/LUpi0CiN9t3nVYuQezZHfrcF2BJ3dqf3Nb33wJyR7HTEVOt5cmdNakPW82wj1
YjwZeiI+owOsyP4SEe98aVmamyqTGDlQFNZyUW0wAsWzon2RpChTNKVRPezt4Zvb2LFeMH1iW/eN
PK/yEziWhSJU+y/oLNlPJo9QJBdzQWC5wfgiB7VURRBEHne9BgjmFiTKrKzPinlrDiyx0efXFv6K
rWtxXv2inRwPjw9HwvkxX/PceF4BiwOyApBrSys44icCC23xVSvwbyDAi6gCrb9HYe/QGYQPmCUi
WoK8FqKHhdQ746S+WlGalqG64nfCnMHq3TWeAZIVJEtcVcfJXhb5F4UsKewcQG9Qn7Ja7o6aKsjj
ajcqwuPQZJCuOTmz1uEHVB9icSamO78h8z0yg7LKeMJoYc8II61QvcpCZGRJ8rARHnueQS3ptlEP
c9cnH2YfZhVV2NwpO9Tybc+ghWext+U3sV2H28Ow3gyK3dbZG+EYZuRlfTRnzuSHLSd0AINlhurb
qveSYJjpxwN1aFVAa5CniP1/uLD8dymvHKTiz76MuH7dq/FoE+G6szeeabv7Qzxg612OZmzMAoKb
8WNJTCQj833/PKwZZpfxgAPblme5uV86anICimk+eB85nVPAF19jV8mxgPN8395LAr3ivP2dnPy8
X9XQz+koumiQ5bKRu7uHoCpWMtMGkxvwmQqA7tICWwiHM43qcNilUcuJ++XKxEwS0/Suyt6PG7vB
t1DzN+Gwvx7H6D2Pg2qmOi7IXS0+USnDPVP5+1iRwDIUhUIoNsjmIvVmWpAKBVsPS1oCk+s3xciJ
3mq1Xeqihcu8IZkrOMzo3w1J5wXDG33PuJKFpfckNLjMey1p3TcNLwc86eNy1W2fWT9ZsI184uRq
rxxgMJ90VQ3se+lUhQyrZVKM2YssgEff+N7ZgHpmGlttSzjxDAHEx4XEER50YCvStviayZm+hIcY
zoCwekTmphtfBk0wntahnRq3XPy5idQEGVT1i4xSqHWh9GcHaA41y6xkgLy2Jr9AdnLhcSyBVX1f
lWz6Wh2ZQ373BRsrA8TmuQrjWK2qmgRvCY7Ct4gThXFG3tilK7YTF/Z5WpAurFKCJyUg5eMgQ/F+
rwjBqLvFG5f4vUtHJTYIWIaSSoOH7nDZbm5vRu5FDI0kyjFyjSXbtSJLZmw8bOP/945TY9PsU/pT
hsqHman/WR6x1bi591jogsnO1wKE1ntVAgVqQRUeSQfzM6hFYWvkVW/eIf5TfCRnJeb3HY12OlcS
2UuiBWg8XH4C9Vr97LQFJPfJYEM//yOpmi+pQmBpGQ0jjNZG473M/O9DzoCkw1XxSiQj689ic2z0
pa9IEWwujRAXy9ipywmQKtPdL/Sv5G3L1kOpCbUhUYlQL6w5vbXjsWKBhjhlpbQLESGd/+3s+I52
iTrYJ74vz2F8Y08rOSUHwgGUFsHse4hfMNvpf4gOryskBt3vbwZDZUzrIt8lflSf+Ez9Q9Fp7GYw
kzz0fSrSirPKNNFb2UIKLgF+BaeNSXg+cwezPn9r8T5Mc+Y4mRkLS+mxw1jznDy1zogwTWivWuiT
c0YQfQST1W9Hzr64B2T63obth+JLgI5GkV0rK+hbKK2I5M9Uj5kLB7nY6wljhgr8SofzeFy3JYxx
A5br/HGrCMOKHWtgCB84x1/tPf736JTo7Vrd8pxx2ib5uc8HWreivEqnz1KWsUV0ROhzcr1gdU8j
fKReAK9dFdikDp8GdHRjKU2eeRg4TeeC8boNedNAvBOJ5kKSqsNaOZRRk2afJjUMtNPVcBaLbpTy
BrQhwdrosXezaKmamM1jIxlO/k6LGp1Xmr59vhx92AT7xZEiIPbVG5RhlljpiPISB7E/e2fhw2o5
rwpSDFdDdIrHk/tdS6RYwRdy+mjmY6JOAk/rwqaJ26fkGM21aXjJ3xgeambhhEEIAyIfRs5/ESTM
5sSadfvyc9IJEdB/LH8C2FAb2k+h2olSxwmoYOpp1We/wD+xYMeZqw0aeF6Aquhdss1zY2oHQgwx
W2d2++iCRBglDs4oPkK+OtdUKpmWFG5FibUiT7jsICwsiDhFSDuWGSVlklJ9l45ylJjieU3f7H7t
JhDnYyzKu7hudK85mv8C6kWEaLo42IOIIrlpziAiNJaHd3zVNvgsCaWBiZeo+VYMgIFTczNiRVZ4
JGIIOwXKV8okGP7l3jwdcSJqQ4yRmqky5vPiJSlR1QS6PoGYNYoKyNff8TnHNSgR583OgItwlT8C
fZNjee5InDFn5ezFqYUpI6N7aLy3bisrH5xJFe8Oqt3U9kl2zel4fw0KTJDDHdbR90x1lX98xe/3
ABkMdPo78oomGVkbDF9aGGVBDbfuWlUJecvLwsR6VYoUtiHphSuniDUkGVM1SesKvAytlnI4yrS+
HV6bd/cAZ43cQq7CNChvGgZc02m/UtmEnxwO1Hvo5j24ZBP9CnlmPLjC/nNijPy3HtgYzKCE7lp/
f9c/HPL7r/lgOYEeveesgzpoOF1576JoaR7BlU5mEyX0Gvimu44sk6U2fi8c2QbYh9w4FtWxVZF6
+l7oL/l8C9hmPkvv3WT4ZItm3SGuZYNP3HnmG9nR7kT+J/jU/JkCzlUwmDiX69kVrAmxLKKC7Q11
fBmSXsuQGMERyc0QipqfgJvH8FsSxZtAwnwu3UxcnHsNdY6nr0nurr4g5Z8E8hx0W0MMlagvrPDO
DpSNJ82dDFj3sfrUm+rCOu/ahVS0icC0RfB7iMv2IqMPoDevrnA7JwzVMYjfMw1GS9OtWj7f8Uo7
corBttsIdrqIpEycK8m/rrpxsGgIpB/ysi1+DMTH9K92NZzzVi0JNWaQSJqA6vwCwUX2k622fOZt
bYHAM+nY38HAUMXdmX06239cLxHxOw7gj/TZhT9YTjmUEOiCGwRot4qYBj7wRJ8k39R9ys9HVCM1
awQ/DbZHsU+1wZ6YxJvReie5NsGUn4kcwzqar6qBpIbxuMjXqffwC8vfm0UUUvmci5kJ13px7Eer
kJXDIQ29gHvGKtX5eJOtMD28fm04H0x0owNY1uuNu00ervt9KZ93foUVzt/jSOnhkG4DpGuhlwKS
jV88sVnR4rxMF0LVGhAxGPphm5GEEkmZHX4zyuibwkOvS2q6aqOjJ58KJLYGRVY86wlkUeaSNqsZ
LZA4DaJg9afWT3x/YO/DHpUNSxEfckUtknXZYRR4V2iau4LEzh7Pa51TlyCW2XBLlxrdxfqx19kR
M8TdLD6zsN8jeV+Qc2UJh/4vLiqYpyXW9HQVDzypy/uvWuipVg/8RTXUCPqPEXka8ZZTKA2VtF/p
VYhzyLid0wnBZ0WkSzXDMv0NI+JAcJ/xW8kV0y2B8NJ9lhuXz28kMnKeJJpJ1K8MrVoruL2QI+In
rYq5GG4rkbzcCtsDAfVeA13hsK8KgMNOQoBTWAbzVSr90/tg5MCjxE2IiZggs3MHvuoXHeYDqWGe
c3rO9Jqep96TSaJ0vJ3EuVBduRIoYM9s2TBo5xmHaAXtMb2pHCioxpUNQbd916cdiDCOt3D4dmwZ
Pk94QHdmq6rxxP61HW42xEv7QutJifRh+ss4U5UONGG7fe/gomdugAJpN3ishskASnftMwwBGa7p
qFqfAXocu1GfcmS4DwELy2PObSnT2t2lw8PdDvncZ/dTtiT0hCqA7DvXrbgOCb819+CS5Ltp913y
kFoIymqHIxEj378eXW4QecNK6oJSnNhABhdQiBK7L4BKkZPBdO3L7Do+dieQOF7TZmqT1QUBJJ5L
eKPyQea/K4SSHp7SWp9Z2GwFEyfxZb9DPpmIntVltC2G/cuKbMZu2zCPKQ5UMPbWY+QqtSWqXThT
QW7KSpwb0LyTwYPdwxZDnQA34pQl+e0AtMWnWhNd2jBSQ/rDvQhnei8W6Kp1eu59yBNOh0LejYyz
8fvLFM+UpRWD7cXUKA9Px7C7EJcbTQigMz6R4VCq3EQ2tXtXjQeq4PUvDmfEJi3dIM9phqgztNAt
eLH8qirlZLJvfYqxpve879DQsof/QjaW+dA1ptV7wPdxjTJ8/dI/NOopz0kNUEePtkoN6ARbRQFP
sGutiBEYD7iKDaCoPqrPzKXGxDAb3jlzplprCS6R5kHtFT0/rW4Y33gjL0Kqvx2Y3/4YHpsEXkhz
sAJljAIdtsrWAFXobxNJBzyv7JywMwy0MDUfCH1mw4mO4dyD+W8D1XDmosRwHq5uceVD+YzAwitE
MZqgcqQgWWC/LfM3PKEgZ8MywzHzYsj4uiH2hrzCGGd0MmmxoNyC/WIO9vFBMUPFCXRAajVtNJ1b
65K4sTjh6Pc2RbQfjBjlU8+Bfv8+ZBgSzFjq/id6pc/TG4iJbd6FDnTI9jrBDgzSUDtVvX9PVW7R
PgXT0oLkFHMrYYuwd2PtdjWmGCz7ZJrF30ZdXSGTDRgBK4Rv7DOHUF1hR+eXeEKZtWdTHs/djYK0
akxJNsaqoN8EJCJs9zKiwINt91y4+2qSJ1onOVj7HQH6T89ukuulz4dBtb4dliFf9TYr+NliSYs1
+yzo+DhsTt2XconBf9dx8oa60Y8Vcx0ie/cVL84DAmTEJw/PvaKB4vfBJAcNliME584Sj0RgPAWr
LNOgqMN4WIpgbWWMQI0JkVUXgiAGJqQewIDPjNEzM5L9AqCZh4tvnXzrKmU0Sr3KGsGsFqf42eRY
j547g2BiLGnKqwA/nVMrj51w6Bk8Wtc65iog9ZNBiRzZQmgnqQKpy4Gbd/C0k4yzZiIxL3KEKfOG
bi71iHIEYArloHx9XADWAE2Uiu4yPlXkg6bJKdYkQhZkqu2zcato33MxP3I3QmYoLlPMkdqKHQG1
mEB3xQBNfVWDl2NrAa8M9dEOVi32ekQVOE0Vp9Irf+ISbr0FKppwcucHADQaUm1n9IZBE7a/lwcp
xbPLCyp0i2QmdKS1Jlks2vTDJ+dedo8O0ES1kjXtH1wt6Sj4qeiW6ElnKHkQbPZwYa3zoy1SK8eu
YDG22JpkegwdWdeTQWUtqh41D/h86s4vMGbjQDFrD/uIthTzOZRoppR0b1lOBP2NwksXeFtwkUOf
zpvdyN8SaevUsznTlxHhaatZGeccTlAj5ph4hEIMRPZjvDDHqlt/vCZraDvOYJD3ZRRAb5YXcYYC
P0sXD04XYVqd42gZhXDpcXTpoDX2jHbRNpUegXVRqpX5pJbFii+n9HZpmYkrwTfAGiol3mu7y0OO
FKeOdvfp9kn0Kd8v4DnmJaQ/optUr/5ePK56FJW1XyaRGnN/s+OjsH11oo4iAbXIuIZJUlye5eJi
aXvmlqAzotTfBnDoO4PQU3IUmYC2xT2QxxlbMFh1mZNewTxiamc3jIcEq0h+TolXCrkg/aRyE9lt
/tR+TqhYlYh7RgzHlonNy4FkuiYBkXaB6VPfqm8mb2ozg8GMvWj7f3RYHE0pALyk6wrkvTFu+GfM
A/yeHj4K3ul2lOE2ZFz28tDZWMaUK2x2clXfAQPnnoDmJ4b4+K6O+54rzKwt7+AY3uPTWsPWbujG
2loa/00lOqRF5mp3inyja1xl65vTDiVxTfwHt8PCI8rJ74mIemneCQcVaWbZooCGrJS8IHQd6tTV
G10jdyFa8C+VkhqXdjbw1A8gT8P1n3NaMX8q2tVZZN+sTbYSXqeaPD69E6IA6lurLEIuqHCuiK2o
r/j0oKa1II0cj9znIe7T0j6YFiDc015uHb/QSRFwasODZO6BJh/myEaCuuMaZSix/IFXZ8E/9BiB
mRRfEdpqo80vlxVkUw9NGwCNPwTbtWaT6snO/J+b1bVGGl0qD+pOk0rkRlIxtbhfQnR9HQWoqt6E
ey0MVPlKQu9ECt0G0I8iNDJzikTuIhDfXXni2M8s4QXt/cbZwJtO41w7G3fgpX2MrewT5A+6rf1q
2MHkZ5aLyqWm9I17nblXy1PDNjlI9Heer1ImA6H1UzNyTYagkDi5/4CLdGKNIp10iQC5WGb1Am3F
K55SXTk5IRHSRput1Kwvs0nVRXSOTUZjqc4D4Zt6h/TQ4K6WRL5MBUuhMwT4iZOP7DHmpXATe+gS
ZIxgQ6q3zPBgPH8eiOoCHffI2je3sALX0TS/n1O1BiK6UkLco+V5BjN4nGlIypLMUsMvx5dSr72N
u6vethIxlPzQI+olJ7SH7XFIXKhplk1QU4khHTVcyxNJXAZ6Pgoa2IvfhiGqx0pjrv/boAejpDZ0
Al2W9/Dhcn33eSRpG3+tXZAB41CHZKvRzsRHZXBSJ4lauPn3wBkuzUVTBAt/65vScojrYwYyNOT6
1k7wpzWaMzGALvfnx3TFJl9bTyEivY8W6mLN5+y5QwymW6U2woTigPQEICTK1ck/KPM6ePCYEDq2
L8mF+e81WQodeiJodHjeEHhNeJzuNfNpRBr6Cv0l1hrdBH9dX4CoRB6CXDbQkZm2+9xzGRwHOM6F
cfp87RWZEQZdzEOPc6obLf3Q+YQhYr+SzYRRL1fNvKePB75hprjtmpSKw1+mD9qFaQSkZ+XKHfa0
plnu+CMcCX436XnAFd3x0qsxompy44sU+OwHJdAMBfBFSd7BOw5FTmGg0sgBzSeOOZfHCjnUvZGX
kehVDmV1pIV/f0Nfart+K6LYO3KUJ8VldmF5na2sWfCPboqtbEUvgG2NHRYBTiNjQU3s4vB8OevD
drjAo4IBVfrNZKcL9SOzSrwuL16fNuxcivaXdZsupBPyanghic0au/On5L6EZeODN4aU0S6hNSCc
vJfMebzXtRB6CEzWt8pUc7S2uOqlyQhEUq1cTgbEUE4MUvUfGkvzkNNjtrrgA7c6cvZyhnnEzT4z
c02cFk84+EK2vVbX5dpfehT69VxiY8pVOX/vpyk33P4PIFjfqJjcnPwYu15R0OqYhTcCKaAGL5Lh
V2NSJAQZK8rDJsebLqPzmNC0Z2XuFYG5mkAayTdSAJf6Xbw1KclG2MasW8yqS7cK4IYNfL2s2Kj6
9X4bE5OYVVxx0ZBtaxKYqUQrUYxDIztobMlSlae2N9omYgUCF6JovQrOyoBjN0TEQGXMhDDdwSRT
82ks6+Z8iZRObhWM11svuYhsdvyK6NBvTQUrW/M1rLfIFp2PW/LLDyDMSI3FR+0CHh2K9w8tddbZ
NMahfBF/MR9cyTwM07zLtua16wyvPzgn+s7L4igHTHggQG+/tgrF9BFGLihI4b4ePYBs8heUeS4G
7+3Ht1yKQadvHk12WdTO60P9YsHaQw3jI7oR3h0Mf0fF7jU+ivF6NuAIseu6XdWnNjbB9hLM5sKu
qgAUka76LnJ4XbohZl8leBCh1qQG2ZdCQO5H/o0hoaWT9JKai3H4pEgQ8rPqnmoAavfSriZKUB8D
90EWmr5CxIJoClPLzuPyxxSjin945inlBHMiXEkgcxYKxOS1UVOg5m+o0Vk0wX710rgQBv/FJtgN
mU1akuss26CD/npyeqFlFbiP8P8yZdTVCbuLoWDWeHInMYzcy6BaYs6Ly+Sr1Tp9eq0greJT7U7n
ce5w51hhE5O1tiZYdGMOxQHS2UInJ4A3K/JBw69A3em5wapfqRj8Qr9W3QGfLfZdiXoFtv3jdr2Q
cQCB6qqqwv/Swss7kPEk6x0eMzqg2iWe2OGfzNs3fDd1xZL/UfhpyjVXWcJ9RpXFQyM02MenbVlZ
YFd+6MGQfYwW4IFNYe//jYk5a6bzpoL5IEZxZZGUm27vlp3ebYSakfkUP8Gi5gdAaU37CH7L4v+Q
0SpT/FnKRkvVXHGR09pIBGYmeQLU8d7hIkE2z18lEhGqG33JZrjCPiYdfKa2RCute4XJQQdzx+Gd
53+XyIKlqMKeZcOFLs08Xh1sdEc0gAZZcdrCwwsklyXeujWnPdXZwHrAUkKLDGRq636cxZ8Y8M4s
HWq/OMNWWFQnl66CCmM3foBj395iMGJyGC36amllQFXMRPIF7Volxv1+nt0FYhPb0mdh/BFqwrFN
ua0EXDdUHoSDnk/YWelo5BC5LN3mf+IWHXK71EZCQGV6PEcycwS7TalYTScui7XExVg92w7jp60J
tp0HvWBTprS0Da2u9qQun9nDOYQKFhMYhgfw9KnPc1V6PiRbNG0qheZYCJviSvjBnGV7/UGwdBp0
C4RJnPE5pECxcKJlEtS8LXCwNmbg9YseBVbYKaJMLgXqWjE96b7yk1rt+Rcaoqwre0HJm3d93Yi1
D93kJsfkGWiFNoG9z0J2KSXkQCFDFTHcASOr8wELmWDQ7eZdfXIbJxZATxG89ovdAchjkLXTGsth
l1nk7xdX5Pwjd2GYqV89Yqah/fRaQWMTYn3y7Fz3doml1x2FEp+Vbt9DfiSnPc45//CUr/732zG0
jWHGwDyz0VxfFjhLDzFu5WQ6aNzlgfqfQ30l1OIc4qcP9ux6cQ7W4EKD36yPCf55TaRvqj9nJK//
QWEBulA0ZT9R1GhHlAZD1+v/MssCt9q2W44XTtkBPN7ANii7/3ow9UIAIaSDQvjFH9TbmDJ9L4V3
8wjwunp8EeBplYzCHCd1QCXH+qbh46RqqLeadPRu/a+ASv/KgBIQ8WY+CK+QMX7JAVesmatMlP4z
1+SOhgtgoRfQYgqOPfsZ9eauUHwdkML0MenW/AK7s5Qcb0awmaMr3zvKdTDBDq9hMgSVSm1QRZ+3
s5QO3zbWPSSVj/eb8P83seUaifmwryu/B9KJzHQGtwcEaH9pbs/178RATXmoRQy7ZZTzHb6rfeKW
SFfvc83U3Nz/1ueUNLQKddDbPesnPMIolHtfQkRnubS1ye3pFMtOoSZJzNMpJXn24uCxIgV02eqM
DPz9TLy+b03LVFYheU7HMP8STsxz83z7iQ/7woH43bFZSuGWzs3X/FcvZ7o9X6/QduIL2PQxEZnP
tsBFpiwg8ytlcq+TAPs9Q7IkPA9+dqQRB8cmHibJMpPDf6uG5sPLFm666nEzKnX1ucM49Euut9g2
ZEdyCDzNVak9KHUgONvnHGNl3hX4xBoT2MaroWKLJxdvmoDvoAf1/wzkGupXjgoz+Anc6nTlez7e
v3m3+sh4tXaLOBFwTkABdbvIKWgz6PjgUzVOQ3D6Kw3a9waF0zcWipzr5cvIQd0Ep7AZh0fJenpQ
VUcMLXZEun4VLtCB20ALIDnpQ/1C4KrJpdGBMyqDCuZl+TAXmkhSZhCHbTAQ5tWBKpU98vLTAUvG
vPekHYqsc1mxySi5GzVzYSS+hAM88nr2jMOsYe1bsQLn3e+jqmG/oE1lsWqfoNMEbNHwTLguXjqa
lkSx6/KHk5A3QCEUnAuwzS/i8BF/JUBRz8XDivavrYed30aWr+TQLed5fUjF9+Cik+aRSYaTCdI4
Q3939drVl80q812CnJBQjolVdeUBwJelhm1HbEhjLKkKwj9TvAdZK/iYqnH+I442nSu90nXzTBZH
sSahSAHQcHhvRkaZ1GFOyNn1fKo3cOdArQ5fVeZEcaECYiRLeL+Ry4SJXTDwvJHO7svuhjH1BxS9
NiSJ45n4XamAHyUPV0ATKna7r42VouvWfvclCKKA+MD0Q3OiPvG+ZazXZwrzPC4XUadzWmzM3BlS
G4jH2QLNnV1+/qsgUr6jHyJFcw1TzspqZ1EwyH4igm/6aZBs6ph6+PHVmpiktD7JM+GsmrWKiCNc
u+UJmjUbwnT2XwjMDfnZ3eXPZ3PfcneZPg8nynzoOSJk6iDzzgpOW/bPz4nQj6z7EsCFzrOqphho
red9SzhyUveE5FRPfVBzKS8N3JfKfG+15w4RrFRXf4+TiLWOCmY2JclOnii+1nCQ2JhIY/7nInHo
i5TlVZOyAbsFZNc+dhIfB7DOPd5SQ5DkR5ssF34ZHS41RbZoVf6pYyMVpPgkE/YOsd+TC1+r1BnU
1SENrq8fPhra0u5L7IjKmZvq/UVIz4aUMn1IiCdxkBg7IYzqAI6BNyRKljWuprjYFX+WA4uMBbbu
7LOlzcvlhGOZ9ysY1FGD0D5xJ9o3/VS1JS5nJBUmkyxD+6NLxzxoFanMBuPBsYialWT3zhGBmbC9
vSsIXVGP6/W0Q66WRGnd2tu1YWD2xY7L8Mn6yC1zdU0LRM1CeEPpg6e4x5e31+rPbYKmu/VF4GP6
NR3hJ7WTacTSDKrqAUXprCwcx8fvIEpAJIoPywsTG1cAOM03FKXNMRliFLR6iLWifnWhB5KhgW+e
ixlW8nNATb76sHBTwdBB9UUlRGzWSkpMDXUxq/pBiifSngA8Ca44XLK+z6dpAw/miXrHu4reRNMZ
FrvYbZB2pGcDLH0uWaLBqeG+QPRHHmtGiQY9q8ieTg3IPWRArjYri/thJ2o2AVfs7kAirlwpV6Q7
GStRc5twUmzfYgegx3EgFv0vueSLZf28NJtQ6gaa0G/hXoSkyeF5eHNWzr5HinIL9LivUIE4aM9h
aEHa9/R0MswXvGeNDv99HAwRC4FS9ESBrdBqyD2nOQp/2CZnTSvdOYM3fNgNgwJW5uSW4OSE3hFA
ov/pB5MVYEScJCSmNCY+KL/rnk12vSglxCJr7lJv6+yJJMqvluzvMelWIG9WjHvh13kY6bBdOdNQ
tgDDJ62ueertide1BaQHYjRH8sR48vnKYkIqMgVTiQWQGIsvPdYvS2IioED4EbositYcpjQH8vyW
D93y03g0IWjmhq4znVzA8gblyVLXelBTP58Ezea0MrqUQZzVDwtbHJ/xhrx3lo8HrwqHkOzlALrU
BTG8S86YeNLqEha6Fy3PjL57XJXbx1op1gG2fm9wHSkvLAdbxygQXQ+n3ZkT0HUdsH9lglKUz8Tz
OqvSKzDSQXIOme4cgo3QI10oF7tc4bzA9TliF334sXCVyzBI1IUwj/FuXUQBv9px4cP5fWsAuIIF
5gAM74+uCSUbesm8wzg2I3RJzKQi05gd5Yjc4N5m2Z/zV5ciF3UM2UovmOg4t5Tn8/2SX71i9aFe
tOrNth9imePBhoviahMsva4yfRhjtYRjq/1mwwZv3CZ5SxtWITN3tkJpi3alAwKwB89H7QORJVrj
QubseqTuShRUvZP1ouL1FDWP19SdbfSMs1gD5feLKj6Wa5roZSuH8+07aJbboe8Eb+dJjglqdyqP
qg5TMhUv5FFtHLT7D5KoCZVsLVZmMODr4wXugNS1LjQBoGGRK8G4DEfVqOccqFwQ5MNI53wDuYi+
G0DtlXtlVJThTCkf/6xbbQeN2SW7r2m9quC7IpkEvNuLzDbw+1SJfhA711NJSblL/upn3CDOey6z
uz2BIJMfYKKBsmt6GdF9gWXU41E8cx48MPV3Q7uhYVbaqXx4wAE+mJ7jWqEcGBYq53e8PJaEHWCA
B6RuODLZJR183D2DTqUx9nu66EF/7kZGl3AWgpZ25+mDtsSrZ8mMe2Y4iid9o0/ejTI+4CKwopDK
Y/FjQyib1jWTpTGvYSgjG58ZuISz1FJE/Lg7rnRfdqW/vtmzcOEASslKdzOFbDOfPIFAvSkakMo9
8gtGd/PSOdU0LwlF/qT0r3dqQ3iBgt5oVnwD9J5fICydB/eR/BiPU8IUVzm6vSsulrV3V7e67kTn
VY0AmWuuaZTisrmW48f45HG+LviTeilrZleB1LL6pvtAGvgVprvQfecBakm1Tta7v8Gdx1pXU25v
V7SJrvuci4kGb5yPkCJtN+KO1uOudQn+4CRw2DARB/9cKh33qncEws1mhAheM77AhTo9pYN9p9MN
bjnp5NUxQL9hnYSWZ0Isip9kA2fibgSUq6zcyAVTIlKWvB6/opRS+RZZKLVmm2xtBZTC2hruZpG+
sLYHLiO322LPTCWM6JZ9COg3TKK7IMAE98yisDo1zEmm0I4HHtLgOu2OIvYup4kBCzGij2rvzhqU
fgaNcuq/IAJvyz7+ZlemRbmU3zC4q7c48D0rtUWh9K+0pnM9R4gf+78om2tg1RDteJ9ponCMMxj+
R2LCIK+xjH4sxnPStiD8Aw6tv2PF8n3R5EyxXD6I/wtb834Oes7ZqPsuK6SqhYwa6sA/WFem6ZFE
CTgPP7aQqQ3TDjXzfddByPTSUaDud2UdoS6/Om35+n0dEOwUa1C/xL4HupkMk5N4ht8WXZj7pCDp
qsdVtKhvcrS9fdvpMYfVm2Svwe3FG4Dv3rt7iBt3KDmysoKYSE5Ao23oEnobKBqYBrwixVZMdjqG
w2XjCjNcC4IOwcyXiM3juXRjcxFUn0Lgt8bwCGB5eZ5LY5DzweQ48I9Yxe3fGxLnMs/EDk9gp41D
og03rAZXD+MKYd+/fYWeULRUZlRibKmwhZ95hqMbD+dHOWl2yJ+mz7Bv0J+GsjQG6erOkfk3f+nw
NZZ4J5ZuaHwqU8t3FSiKMIprXsAopiG9YRBDbOOKBbmB0lJg7lUYgaNPj56u8i3H0PYTc3saHmMO
pICv3f6vWjyYCjqk7EXC9gve8vAGXpy8/tJULicyy0X4JraVM4eMJqD6pcKc2jKpD2/sOmy2gE2E
KiMKSehMc2XQ+VXlTcPPzN13VP3K2NPRX+MCdjn0yfjODI/x9DOCPUx03cqwEsaWl75Kh2NHoX8n
0BvOOm9IntC3XpctnuT/seP875x8U7NTKa6YfjiNTh65szp2y+k+KsYUdYgiXnUO4GBkTtdtmPxG
HSu0awV12VsVsMrld9rPJklJn3SnR/e3u8lCZDeMh3TXcIaOmIV7KpSyL2cVj1L5ZkB2CQxL6NO5
MAfwy8yKLE/r3K2aGlT42rrb3jyi9TjaJjRGkzouijmaK/P2NzO64S2Zlb9RwoJjmoqm6s205HE0
yu2n5lIfl/aqPP6/fqM4iVyOZLGpScuzJIXwpwgcD1jgYLnx/9IlzgLG/0gIg8G4OOyX2xtdlC4n
UCKt4D8kisTplu+uSuhZJx4dUUetU1h2tt/vSUAcq3BD12S1qWmD7Y5tgAA15K7LBeEQ0WlhF1c+
RKs+qRG82ewNmVAKIsL49ZriiixIODfqFlJ87VrXfUXoj9vcV1nvOdGL3kQogZyL2FSlBhUlKLun
nYtKJM8b64vtEsNUSbhXw/ezeFh8abnC7N14LfmkC67quPFna4VbX4nwBk6meZHxpTTyT45JQyXG
bVwuUhAZA3JD6bJBMSXYt2dm4F7O1cq0TRLEM8FrQb38t1edj2PLiKlwd6UqbS4VzukBLSMPgWld
qCMRdD7nBHst4Jt4efJ/wo3iEDI6oqD/eAdLs0jdfxRQ2aWNpUowA69VEHgOUifHAZ4QtTZJZP1C
+IHJE52wtNbWqyjyOMtP94TWSyyxcvlyn4wt3xgB8HOxutGndCOaroDH10DwWw/9RUzaAKg0edmU
qoLI6RHc8+6RqIdn9v3Qjns34V2K5uYEF2NOawSesz0SPrs0+PeToaVyBH5W7KcayxQsU/Qs6/nW
8L5wgh8hFuIxUlYELJiWaSvOlHffs9ec17hMy6g5teU54g6S1dr8Hg87Z644ezFwygKKK6O6L7bT
/kvohoUzr+lJ6T1oZRB5aWt3Mt7hw4VFwi8OeM+XrWS44yXTmRiH9oao5oJny5cm8C0sACYN+hDJ
l5xO3sR/TVS9jBG/Qk5h22kdYMaq3uXHB4Dp8xX6uF0H4WZk+w/dY/dvCECIaw2C6uKlfUcWMqLN
efur2kSRlf7pC1z//NnP5Xwp9wnkyP9GUwkUfKdtPt5t/mxqIppUUGLsiZXS/OnhBS9lQzS4JJ0W
kT41mlOBN2AhqDmP4rgb58DYTAsnVUbwh8uk0prWyn3p6ae2fYO3so8QAhKwAr17YvvlV6oHSYVl
FBfbGSTjNLPg3xXFK8QuPueRQpuG8+f++V5/PEdvhqh6SnMpFogQihtld0HCjcUiI1JxYLFyrk7G
ZMGZPIJLYHUhdBOdfxJ1L2KEvjyG0oz78n/PbBh+KHkyTiUpnB4dikggJWahDyaknS0fLwrZO5+E
TARTWn5OPbzM0HUFola+GWuiA4WKfUZbE5P+Ye4W1DXDQdcjtwnsMJXOe0G4/Tt2NBgmkiyGugGc
wnbYgZ4jf8bXUG3SYb5NY5wZ4xtE1VHcSMPruoSaZWMrNQvSnT6h6we2vcgj0fr7EtJPjRv2CkxC
qwvxptgUhFLcpmT3puEM2CwphosKnEK3qPbqUtAS+AF4BiBKGu6NU/jveH+ZHynrVOh4gwmcB251
5ddqCUUt0Mc91fPgx2AQED3r3nMk7czOJJQD6B/f9WoKbjXtKqHN1CYxnGc/QWXArG2w9qWwtOAf
+FrUfGwBCrc8OkccKJjwEt2qR/je4da9AZjaMW98WhHuLWlCeTnkAT4jPDxw/xwoTQnMXPh4eFAu
ifQZH/gK7Bx5H4tpD/seNoqGc6G4W0eb8qhl2/tAUn9H6TYTreCTWLYMyUEsNBNf/PQAKn2v3RT/
9msrCmY7UXPgk75Sx5mwEUhfudv5FDns232ev2MaOAzZZ+gs91vRdz+l2xBvdRO/BHl/y2CzL1Ef
+0hAYu004c59vf0buJNvFZyxxxXXfieNGcHd+oGLB6y3mTJPFcM1u8XRE534J5FD6/hHW7DMmfUp
hpSpERVsmGQVEZpXcsbUkS7BM8sVT92MRi8VoeIRhORTOKvtOemL2TuSurHhXxpgEM7XSrltxsPZ
X7IDU8RdXPfHvh4J1uNA2h+LyBaF3yAhMi3TFQsijGkGgymA01mlfH7KHktQ8hH5lcakuFSWAcjy
QwgBCk0FgmMiZIrJ3hYd3ik9dttfg4ytJ99dhKuM0iciZCZ4ainPJEHUFhAcJ7p8PWiRgTXE4q4j
LOWPpntFDvsTf/4whv0R8BFRPlESUF602JhLK1hv/F/2r/M/5uQb2Yu6kRxO3qgL8gZI75/xFNxW
dLq8S6LyTUPGN1yA+iEPTSEebt0KZNBwU/sUbyOojKAhKeKVmdXkZGq+jHuFxQzk6rpb5/xdIqWO
VQBAxYhLxV/0zUjUsIap2JqVyIaKTiycYqIc7BLy7gfEtmAkQ+MGvKLto3EN6zux43P4xNij6jZP
GQA/RvL+9JxoxvEELnXMrWz57kP/kYPsrzLGtRePg/pj328v1wtYgMuqApcDAgmVxKfsMB3octGW
Qhf5CnfzokHmX5NFnVGuTF4ChGmZ2bRbGTCgspOTNqQlmlFnjrH/GfNJ3kWoBREgYJJIcgFwzd8A
nfnVj1zU2336QXPbRzhbwg6twdZdghrld+RS0MmzKrIYthKaXFc1xPPCY4csy9oLc5DE5Dbo+I/1
kUMr0VkbBYImx5C5HFt2N7SFz8KA+xenVtMlRdJnb1XzOyUl/OBhYw2A4k+3a0ZljHecgJAGObec
fXx9eL3P8/CXbexAGsr6VAKh9xVHWKq25IHOHRBhZKwg46c3kgH1JMPmZt5dkkI2p+bNQ14ysDp4
xjNLuxk7unZxE+qi2kEMMaamCcG5WAvBymHhTdAnslCYJZZbXUHvSkmyg67weK9ZyjP7g2Ij3DGE
Ut9w842zI6h2XHwFj6UPAd1DRZ1K6kLhwFED3F3uEwRRUc5azuomma4UPa0+e6vKdqilU8uX9dde
626DNdcQ1yVi4sAcEcX5HUfdxRry8EyL0jL/3AQi3wOm6BCdwOf2ZLJKkC/fehtMVh6pIs457ri/
zH2f60bRpYQ+oI/JgjyFAearQPac1/JmmmhQyuPLs4rsLh1Y9edGWxVJNLKzyxpusaYZE4bOhBsV
btv8QOyKtCZAi320xPa/zOHAYyAYAeyjMSx5404rKByXrbj8zQKr59kJPaaie4ukbypb6yPFImzf
t7ca21oNj61v0yrlZxNP8gstSwslyUTqWyD2J8tM+aCtzpwfAfV+GMS9/AnsOhJ7xcfCkW4J9z5o
Pgme+6MNCmmbBZU0Q+P+r4uHhABgoN6Z1RckXZ6y90zXWhPWRCmOC1bFw2fLrTpWpoCA8alolVjP
D6kVwgGttmQA8rl5uMa0oEvDSyMXRW/yS8zkVsfUF514Iu3QUzOCD/4Bkn9cQZ8YQBbOIt350Yo4
oK1lCqm/vYNdJmFX3yTh+dGNiH05KKk6MoERswYfsg6iBzXRbvu5C4u/0mUIcI5AxYUp8inY3xXz
v91yUL3RcROeIj/wUDuhS6Wo0IVehJDgiW+ayly6LtXVfVa6TSJZhXsEo08sC9WqlWadM33Ty5d1
gqup8aL0wNVrAUE1z/jG8aKs9wWak6ayynHakh8ZD4KfgN3MyaXUqjuZhcrjBSb73PI+/2XuZV1Y
8cFNZv6CTso1UZJC5tXdkEKC5pN1eO83jgfXWkSccgCBeRkjgGDDOfBW+Mb32s3/Ims+bhuLc3QA
KWRL6RAZQOjU1zEfc40fmw7MRXkRxdzfySJRBqjMjBcJrulPfzYAjELlDtrrITuWIvp3vTJuPGlK
pyFHQEqXvJUEdbrtunyxXWBXK+xyTEFDYPVXmfc0vRcGc9WUDACkEbTYjZZAeCRvYeCMEGQUfiEB
JLl4x8zXKdEOyBKs6BN0Dxn7wKrDgLNuuOvjRvIL/N97P5sX7QYFRu/h0I3FNtCYFbFoq/phYLWQ
Z35SYaPaZSDPYFQ+GwufGdyAW7HwyjDmdY6ULyBvzzihh/msyhKZWz8AEjxWfRyyYC9qXp/VbtHv
CY8Wu0R3biXM95AkURwfBqwVVcp0EzKWs/sNyZFjCh5e1cXxHNhNhoy91lGG84rhllUwjTZHGG8E
b8SVJv9bVcMRYJtxKP+w4kCt1B7H4WTCC79Dt1DEzWdySMi1QY/Ex+1GWO2UCh/HU7xMBREtfS4i
fY4j9KFKobFq6ofwk1J6/UZI5GCrC9WpvX+bh/M6nCo0TRPv8uRlc9ZnfjDf8J0MUonj0gcdq4eU
4Nz8uYNVLGlS5MwwuiJ12AuaZmgz+H642G++bDzN5cSGNO8LgOBLpM8m/rnNNnonAsKiW3QZobGW
MGaMfSeFwROltnVOIK8ZgKIHF5LrHBJ3E4myI9ur7kfpLJMajY+ryaaX0J9Ripot8pVZxAaa+clQ
IXXMzCe/MDzjtnyV3brfEedFJYaQCxSzVxALGDdP2Z1jtRnm8+ixKk8lR3ijVTxJe/sopoBZUbEg
gPkHTpGYAyrEfNIDre6bOaioK3HB8yiiHfkN/Uq27RQrHcXc9r6ijYc/p5bnJk2aH+L3t3zGGc7h
1+mRm/5TpmWNb9f9H8V0Z6WU+HZe98W1ilUNE+o2SPVkIjE8y6VJejyGmKKAEKDDujnO9WY3oVDd
W2YqVWI5xf6cGjtxFRJqjTpA4e9CebpCDhoOhlS1LBlp+gHmpeFTK5rplPKkPDqnoC0dDAMikU2l
Id9UWsaAOWESKSD/ExG+LI0Ub8xMVB5kalxiny/iFYMeB/DlUPHRz4J3mRIzty3LojRpZp7I+JY+
2htcf7Hw5k5SFRLshJ/Q3FjoY0PAYcz0rMwBxdYMk4Ow2AiNI+LgYVttwivfXInEK5igCK2mha+f
+QEhwnoNcfTvAqAEVKAierp8nhu1O4QRR9wYxWGTiUpcU+s7X9IlHqQhNMW/ZvGmKEvvpXhYKqJe
JO4kjQWpZGZR58DHtRwAU95FhyrYI8sCE9l6vOcMSb0HYP7StsLI8nt4rEFzWWjmW1O9I6t5pIsu
BOIIMDs4DLRF2Tt6Tu3zSy3liCXvbaYU3Ml1NVwaZ34yFoen43tm/I7yb9S3BygUdFvyEkCutPnw
lrQXYswV2nu0xeSiZ6avt5URrxs9AqLlHARj4+iBnAurpXziHgB2khr3T45YEPSTJ7EZObHY1kPs
IygC4a9ii1kIW+9mtNINIhoIzPSCpeiPlgdqfxot4LBrJMXVzjhET2j1waKRptcoEvN4P3P6coXs
uOAKiDpQz0/fqLkBwh1mcwJ0HgbD9fFZslSl/a2jAqeVV6mi3u+VJPMzQSuSFQB2Rv84/GJci3mT
pblI4MAabxk7Z1OJ2dNczk6lU7U6L4kYi6nUJ/K+GFT4DS5VRQQwbHo+cn28d5kozVjmhpXSdNhh
uvDO3Kz2MMkrq+bKDIulp5r4Bbk9OiBP5cLxJGvKmp7oxg6vHfRgpeQLGJNHDsvYGiCPatjh/CV2
YmClzlmBcOWVn5coMyXfEvWCtPmLj7/Hhnz7LY7De2p07zJGGvMyyTZadjequWenjXB6qyaPOBVE
gRqzd4/eB7EPfhsIN+cm0Np5fBXjog5gqpCEIoK7FmRCGz8RkkFlUaTiyxfXuB6QtggfpsrrF9g8
ugacjzDBkTw8w7tR4GuYXH5Ny+UYTptlItZu6pVIiVbhYXuKUgNmxJxNvJUvpyMTdm7oaF07Kqm1
xdkzTokmWKWINa2oYW8atSwg6Cbm3e38JF5hgtsTG+oRj3NnK9RYPMgknySk6sgOHUNPg0U+/6jY
GYou+/OkS+fSCf6GoLR+5EPN5GcIQTcN8KAXTF7CuPv+K3gBVrqLSbd7RJcSg/keeOrmT9xiXl2N
/9FLVUwgxeLs4zmHMyqo4XVo0fHeO2/nWFJBJEWq4qPm/8OH09l09ECpn5cqgkRqFrJa1AUuEvbE
T120g0IlWWH7DWfu1W/PSg8+CWm03V14gKt+CPDu/3YsYdvfwrx1hMXBCSnE74y74ew5MSjQfaAQ
cLFgItVUGtSC9GnUohqjs1FPsxHXKEp7jvEdNZ3wThbOWFjYKjFvq4tyCZgd0Q7G1pwDDIbnQ0A4
PaTCv2/g3xkAVbbSIUGJyBR+jZuH291W2ezshpZqlB5cjU8hzbhTwLMbV8wD8ENyM/UFbP3lkvra
ist0EnXdKMUVw3fEzZBcZO3Jp1zl/dBH1XZthG8j3bUuq/NCct59ZuAMVJhVh9HSNktDYG8loiqC
Yxu8bkJ7rg+3yZ6VuGTsyw6PnqDCDFZgvtPlwt3TMt2mmIVmNIeS/yfGfvDbGQwxgVln0cC3eH67
Djk8ZqfS2NP8dSRRxCmwMjDmBH6uBi0ol+oETQkN6IqjvufKpO1pPa/pnhamkiEDu+GevvN26ey1
aIsEMD346KBN8lPo9+FId8zImki3KKhEkuwyB7RtkRBnKUri7cxkIXcJK0J5JukANnIONsu2V0mM
tORPnMowZWZRrzrDkzeOBejTqXzrJ7aMxhn8G3pxxcDMj4b3LRhHRZcqZoFRbL17FiL+bTv34LHx
2gr0KgYafRFH7/pCch/m/sf3i7K0bfaeVsk9Y1be/rj6h3iPfQQiW9Qu0T0w6zs3qqd3LrnckKTU
QaUr5l6QNCjBVYjMmkdAZ8TfpAukLdFBoZo+g2tSCHNq/jtTrdxHwXwRRZLjUNvVFL5gqbGdRFoR
pjcyw5fw8UlWTIoxVljUmcUqwXYya9SkbdzPR/q81VjxsS/eJEGaoe71+N9v3zNGnNwJPKwjcq6Q
s3xJU7AFvE1Dy4+iC7H4MyzwwyzKlg4IvnJBgPgtkETJfKKdIbrEAVv29nymrJwF/mdVoj6e1Dzp
caoBFu4McAXx7YII18pVN8tPjkhBp4gtdJ/Ir0OjXhLqGQK2nND7Myvs5tjOU67bNuDmDbf0WK3I
XbsEh/T2kwnRJvNfeMN1TAx3VKF+TUXSitdL/ZkvMU85roF9y2HBo38EWF/47vl1wYhX5wU4jUrM
CZEK1gYCyB8TTYtE1jpNyflTpppoCNT17TZkkq1+r8esAwhIWC7pLchjDId9t8tx4cNKdiltidLt
UnynyJAorKvYZKG+EhUBpCSRjyaQDK8fqaCkvcOLUyGNduXOspLlaUW9bwBy7G2HJhY79+TE7u47
YLv5zDkrpfhdBlSj/+9N4kksjVcLS1LfMgwexibf/UgBFVk/HTET959DtbhdSUTvZ/FfJWIuqdri
SCYJFo//JOO7l7bbzAaOEKk7CuIYaTTDhROp4i3yRm7VLCeIfi+kc6iiFg6VbSBmBoLoMhypY5Y2
phYokcxtKKdB4a3XEhDimcfnEQqslrTFjTJrMxsTrj27VChY0tC5/CDSofwBYoC3IJaqdSnsYQL6
bOFHuRfzbXv0/xeOH3VuEqYaVZCJ58boQ4F/dyc8dLCHEHhfB+3OMW1R7NW7Oh9FJ0lLnrP3uZFF
bg6GK1XcKc8wWr+mSLP4vur6APvGuOBwWqDv1vlhq2rSLrkKKYqX/DnKBRxNj6rIHAQPk1VbDgNw
I19BHaeoo2YCse4nCms/uBy5eBtX/5qmMsgaYuH4zSNZstw5ZXAYuLJQC7QbTbWMZ4mECew1CBwo
dd7/RbdgtNQDzEaTgPihkuH9ZiPbxXcIJ28CMKNie6u0Tr+4/fZrZmmm+jQcTZkRDCos3Q4tmfo+
Xu7Q5GkkS3xBJmWOb6tSbfgrCkWv6P/ScPfInWv1XAeSTXeXqz1HMpyp3YOtYOQJZeGiE+5x1Cuh
5X8Tef90eK+0JXTmMjKt4yHjP0CAM1PRRWIIEgT5cHkhBTSx7jUKWj6AiRkoMC1RlQPg/vT/V7Bt
Gw/ww+6cxheWgodYMBXElLJUjOjroD24TXMUwwrZjE5+2hqkRpeL+eUCQR4EozASxVIFXAMSqV+Z
7cuLR9GFAnImswjUe0QrUFqC9yRnEB05GLcU2jqN3wr602GSSf0CqP61UZUTD+8uVyWDQK5nUBIf
OHr9biOlTQZ0TZ4OnfakbcJLqZzfWkNC2VceoHsu68V50qRMZATOeSzofNm0n5Epz/kL5PM+j6o3
dEBLySiinblkeNaUoqzrPCR1MyblgLMEfEVI+So/ZjJyB9wV9KF579B9yo7lQG/YjWNwylcreejl
tJmjyRa6NfDvu2RgGollbt3pVBcE959xps/PHgF4IFigMYwF6/3nRd1wHYIfwvSfVEC8ErRxgODa
wjRLdjRoBswJVMGR/hexwsXSoPyjMqVXUUf4WsUGcRn2T9AzP7/nTZ9NtYBDHI6dgxFe0fgG20sk
bMrHnBEh5hdwqEMq4aaUBdvg6+1gIfo+gNIQmAn+Gu0LBkuYMKP0LDFQ204DUS7B1fU3ci3jz3qn
4zTQ+Dcog/VDga6JYcmLQeISf/s0j8+yPCaRkULg8YM43Jw4Cx6f8rshpvFszWIBg4YoVCd06P5c
mYTT8Kb4jdnjR8Xd0/qUqBKLrWu4/VZttDSVQMeRVzEU78gy82fh33I+llRzIhJwhR7ZWJSn/Idp
HUttuu045dQjdBNYV9Y6GEHz4CspTUWZDj8CV3R2TVHoGCEQSG420DcF/0W3yk1gkFPBBsabr0TY
zg/3uDy+EEuQRFzAGfK6eweUkZHGsVBrTzwdF90XxC2tsecHAYraxt2S/nWIkqAGxF1Ofa1nHM3k
as8udwZ1slDozetwDQOw5t6+RIZ1qYiRWgsLy6lmYct2sNIgQ26GZyB7nwid6t6HH4zXyFjNZWNt
PFrfPrhNRekxL75IW9Ledh9L4+vBXaiErpeSzCMc6T/jNVhEkec/etBBgdrraNcQFhFj+QAZVxEX
MAO5v7VgziiDsr6OdS6AytrMEbojd7/AiuMDxhrQiAgKGjlni3ZD+hcQe47yJWgNeWGSMq3I5pNZ
UOBwmkevVc8TLaSiamhZyYFzWUKxcVNtGi3DKc2dv9rUORkJRJYsyxYLJvhFzxXcdg2WaOTyLrgp
U7FnLCy1RnWqyoT6WAX4de9blV8OK8lLWCPASghsQvjqwX4hofLXxrv1j8aIEyconCDiLutXkeIw
Ys+bmNrJPJG68ZV7dUL3GaQqnQn9gfSuEOAylM28FdISX9aYeqqdm5CAB+quSItOoVROtk1/tkTU
J8k0XFV53ddjOwznxxdm+yxQ859c4KqXMOZResyIGXwNdERR30Fk3DBhiyaZaBS+7FgFbL1PyviA
x0QfVxjs6m3JkKnP56Tz9FURWd3LNy+AblX/MgQMZ6PtELs1BHYPZTqbqCP8/FDqWGjr7CJqsZ3x
bMNt3+N5KBEageVuTgNWxcSFqBIKlW/5fl4aYPFH6FO7Ap+hx17pen6oekAd5Odb0GiSN2hHXiiz
InISpNO1fWiriRpesB0WF60b3UzasVM/xSVhxV5a65qb0gQ5UEwRFN4lluAHH4wkOhUTo14RovQc
cD1SfRrrvcyPVB4v0sVsH7dnkeYKO/dSmwOSuubmnNAaEfxRs5rLL2zINWZbp1f5m/wHpGN/Lz/q
/wzkEACdQN6Ff9ERKLL4pZ0+e236Jl61r1MCIQ0iXGFW2tx57WifLB2GhZcXAo+qL9yneMwZa2Xe
QGu2/ae5MGofgdLj1t3ZNEIq3LtTvfLK+8kJx9eA0z1MOr2NhkMhw9ZcFInwFmztx3sx+963bdbH
FhpMOQjC47do4YbFhFuyzh+XSoY7RetNt2e/5uLY67s2NLrlZVMIX/84225ugWiViclZt/mbrTyy
8f02W2Zl5MnugLkcvuqw+UcxDmXWbu2MVB84GF/UMKJsUHN/cdI9/hZ53METGOXO8vjlSj7jUffh
iSc3Xc3j8TFRc2WNuSd0kvNNUzJw0vyWARHK5hpcCL5+DVmyV13jfBTwOLZ67UWy2z0sLmynn1FH
mbW7gFG71Jaub07aMoUjdjtUn78BxC3rtiAC2y+Z5hX7iSfiCOdAq2RQv5XSidntru3zUrtSBPVi
niOf1NA82eIKgHSdxzNBdG4UVN1tJYHatP+0tt/S7IVkOlaFWhA3GxHw4fcRwyJENXfgMF7kPVr0
CiP0mIKdzeVm5kApbci+AdYfm8eqf4hNCNZfJuO1jCiA15byvtrGrbgWrFV6IYkuk4WyWxVlfHYb
O+P7/LhkCQznIWvxKCcEKNoBA07zzoY0PF0z8JhpzGt6xuAyZAReuqknB2r/btZDDrUjdprIdR4/
jdodMZkjS9ChMDqjZPPlNxBWK1q3o9xRcH7UtOj5NG18Ub6CaI+U+bNkpz/RUrf/uC1WbgV4Coo1
DB8tX+HeZ43WzgeLFyeVr9zsw9M8F8r1Op2GZQHEVLOs6Pmh92CTkcNwF8iqjGOySwMc6RFotC5v
zgjexeRALXZK7P8yalPJg1kOgIp9E/TwjY8t6ilK9zmqgaid7FPUw1YPKufbmRni/E+pvG12GfSR
ofMesvMPbp6HrnZVZAj+sLN58BRhVW2BjyLKBgMeEaj3D5F3cGJKqR8PDHgC/IB+ZR0/nTSBI6PR
S2F9iklSLVY5oUoVwG/7ofHuTs4FzJHM4qsMfbiOJ22WNapNjERMLIRgnpKCiugtulHqVNiZRlr2
kpIYCSkGbguF6pRn1Kk9BpvNY6YpQmgzZz0nWxX/uxBtD9CPZoIqKL2lH1kj4uN/sYigxhdFPIFy
/7Nh+ADfGJOwzz4JtDyWY6sX5/11tRre3xHqrLHDbIjHv7niih4wAF89jj0nbCqUxPC+RJCheK3b
yARws9jov/HLUfOOG0Z16ALuduEVPHfowgKpmpe4uvIdqmaCZux/5JIqfu2ljH6HVM5RtIXfI3Cj
/fsk2TsTYHDpvHRTTwXtbeN/71WUzrDSw6q2V0NOeCWo8mlKd0AYqKB4nrfHYE+FSLOXSUlYfuWU
62XQKO+4EYhUfhHMRRZWQ55thKFoWTQHzvOxLOALGbAl+hAexdctiVu0uCJv/82ydprnc/K4ltPs
BWOxHtXgDTN7uWV6tuKZcs/ybuI3Z9nRkC6ShD2t8fzRdU9RNN4SAAKuMu/3WehQwHMP8yNlX19/
0wZbWcoWx0Iasoyk8Hf81i0g0YxcW9DldY91q3UEVQNgnxyzR++PFAuZ7UiuvjxwtOyjy0WR4qfE
NPqT54+NCTt5qRMOAanH6Ri5UN5H8cyP8/3HVKhK0ClHb6AHL4mBAvHJ+ya34PsjLUcQQ32sU9df
SsZaBJdmSbOkvOwruCcSV6d+XfMT1RsrXIN6eZcE5EaSkXSDGJ0f6OCOOnvosxsF0z0chyL+JtAZ
rENQbjBzTnSmw+1PSgoI6GOhjV7TJkS+CRUZzxKr/geC0E6KxA1yfLsq58AC9zkQdmMS/GvGIiY9
k8+mBXcti6FXR99AxBXL9HP5iyFEgzUax4R3pH+V/WaHMVIJwMiUt3jtZ6ynd3jlakyIKPc9T2gK
2s5tiC9X11pjeqWuPreeG+rEWzJRdszv9QbrJISx1m2posIXqC0YP6f5jPMpzJp1w4y6jnGex2OU
jwgzkNAfj/xJgyeSKgS2Ryi51zopISxDsI0/Msf87n5lLf566lUWnj+2sHIZeOmoT5a7uGBJrUKi
vBxZgrecrK9lIOUGHDY6Jl5TFLrlebUpVa261BU5fp/73VHjTlHg8pfP9jjAZPTBo4uLH56PogHY
fNLI0W0yyVCjQVys5DoBVUzPe2Ht+ZCh+rpK1tdpMKVqnXJEai9frJ4epd2kHr2cjCVcmg7WpbjZ
fzI92STsDWDoTNF7d76KwsUJju4Tw466R8MuzBD9RvMY0n3NdHUVBXh/By9Pc6LsH1tC5FQcOMjs
u8mn8pNdW7gyo/i5A7Ul04/6YJctNLvgcljJ4dsr12dftidASIUWOzdZdNZOVVd7kgjJ13O3jft8
tW7CCPDCdLE+22tgrjmyZGudRBh68hb5nLHFvwathMkR28UGPMxLN5b31CzLgrVu3+dLIQmnDxVy
ynXdStCFs/dcnJCaiBsyfGeNfxT55uj171hZJZxe3Vul+X7Osb4LM3re6elmx+ac08JYoA2+Zo/o
cfwjfmjFsCSe6P3S/bIwZ1HCmT8gxIz705joUxYQPt+OQUndzOKEbCl126ohgRI7kEOL0iD65reZ
J6KPwkXUsof4ot+2vzB/xvE1c9WY5j2M27ma6CiT2vHuJk1j+nCcQ8C0yuu1EduNsRlgAewLZxC6
soHCSCp1oNn0xqa/OQzeUjqMZ4xci9RcIfewGpE3v30RUXESJL21gnZtMQXHzf9kBKZi0h6BlHwR
UN2edYLDh63K2oqt41M8CFAmTVZAabq52xF6M1jCRmUY65kViUG2ceUwzDudY9PXevvWHyJ0kKiK
HouxUfoUF7A9KgFU0nHzHNBGvNyHCReLCuBdaueOjnAqKnAjWi2sfevYdGX+eJKgj0Qp5NulNJnn
CLBpLkOuhcVH7KTXi8oI5RfTiJa7ggZLRdzgvc4+SEK2MAapDs1M5cuHvj43+cV6gFnpDU+PC6Z5
tJP25K2AbgT+3h1cqy4/EahNqdt+h6KzRpEIqLn0MUl+f8yg3Ab08/MTWQYhHDlZXUE82+v+YVRv
xfmwpXr6YN3m8EJ9rF8tGD4BRpEN6MR5YQtXfYJG7X6nAgVsqkI4spW+cbYA1QojqbWFyzOv9Bbw
NNx1Sgkes7s+XF8glZ5yR7Z+2sUlPmidAEA5lswXqd115La5T7ILOGmIAxfWS/ET6VoasQrEcFj4
Dctj9i866aP0ryhpvwg8xmF/9OcK9bjGCZpEL5wut+PRVqbRVATGbvJe7jUKCpWJYL3m7ptYU5GC
2lK4QnRR4gdH0UL5o9KCGf01I1RzY0Df88O7C1K9ThOj8flrd70kSzcox3NNBcsMWxm5pn/qB0OR
rCLdiHN/H7bcdYpjggS7v+8EMAVsfZRzx5MB9TJ73xg4q7cNp6gLgHnHlCH8RmjiZcZ0NmAAqHXI
dfzITFAU3a8uv3bc5caWXcQQv0GbbU/g/inSpQcr/VUesAZUTVh1i4PUxrUW4WhzfomeE8rifbbj
mbnph/fU2iimcul6b2bn3AaHIg92PgqSIKkcBqxwPES91LM2VLhjrSQ4SmelEgCxC1XPR60mb18p
6KGjknc+VSJ4pYaBJpl9sWF7tO2F/tAVDwE/BiVUQFf33DRssLhpg/cxxMwS4A6uZOTb4tDPCYfC
+v/pDCbWsk+bXR5zbDVJBDe1O8R8FI8u/ZYy96nLE7VzaLW7yGg3ZUF12r3TwfjfPjB35XuvuYK5
VaCqK/CoqzV4pKHtS3CxWAwxyycdfhFlTSPT/pAvcnLMqKvV4KiIjIseLxo6PzM5o86VXDKpyqgr
zuv/pV50D6CuEbFcDf4ZXy0LdSQj7LF4NZLLBlai5kEPeTCAmMhh1vAX+mhBWtmZ3GN2ybiYXZjf
tmM4+4IPk/0UWoxMg0DWnqBV7vTXpS9itzDiZMjMbvNSyvsl4b2UqR3rgyME6s9cilZLoRZyS7yR
xWePROfn0WfcmxQj0WWTgxGE0N58tKpXApDgW4943woVUPYhcNJb2Hs7tTaRz8M91wVd7FE0P2qf
qT/P1HCHLu5w/D+S3MbvjgElNivelzM5fKrZBdIbmcEg5JuC/DfthqLuV7QYRYUqBruQC5ZYlP74
VzHh6Ynn41YWFquiao4rkHP6o/HOX6BNngty43oygK9jpiqI2KyopbsCI4eXIbf3HqOganUg2r1m
glxQImsZQkde3I5+LUYa9V7mIf4qxgblmgDu0segpsreYyrjBW1aGfmYgWYtHEl+s5g48kJomrl5
MCpaE+H8cVNz6RfaEfIAXsjjZgNjR7Ck3A9zuNmeFDEqsLyQnGmeb71jGzR/APsD7on8GRhU8SEr
VfiYtIkafud8Oc30Mc/vindpKZncSbFatMcsOxR0PpcZRkXMjgejOR8nIPYgftk/zwB1ulSeHk1j
hmQmV6VAjGJrJGikGD8xILkNuvB2aeEKZ/wZCt9h9dmATFMMgv19dcFQCjfxOP2/k9KquTLAGDjh
6CboAyseaXX+vzPK2owSlBdodhZU5QnZ8nlML1vlUZdkFPEUy6bA3mHdMfJkUlnu28CHpYpshnzD
Lz2BPtpD/FbeT759B99C/lxfrSEnOYvg9OOPjl+nkwaJzx5tiJHctk5+lXuHDfJKzRxBv23oEpAX
X8yOdODdPu8U3p43+V9F8G0Z3hpwAUNpZmSmyNjBNW62LPBvz2gksDrlzy3VXv79l6ihzQEyVhDp
SQnatoh+ftAG5WrifAndPN0L1nLLLpdCOCh3wyXmwTozx0GFadhPOtCGVzWRBy5l4vEh3r+HLelO
8qJAH8d99PQ8xYG6v7RyrdmMJwNUCZsXhQ+bOoWrDs3VuenhmBls6WHx4eGQQc9CK10OTPclDWAL
smmHJ5cNqQfFJb+31G2AUaYXIpxUdBscg4/xmJwcixzpqhwRgUlO52yiNDpAGySAYUGINu+kxVho
Te9JmmABlFC/14WcD+PVPo1+66MDk7yjjrmBpd1CaRXncso8BcrlMr+0xzz73x452DhB0sZnz79Z
Blwg9DK0xgtUpq4tCZVH+yRZmZcZwwPbomupY7rCZibRfFy+b2Rg8bpgx5ikfw4x1RI5x2Uk69ly
D8qGc2lrkss5oBJmVPnVV2f5/sLbL1Jj/U47hoZUinyifCsqcvKNlS1ssjM13qndRJwcF6RloooB
5rXQ67876LgzNNwRN/r1reohc/SP/VdSSAISjFa2X0S7ZUUYNV+dfRpCcw6LOgcH4XYKYU5FiYqy
sD1iRekvMJbqMZ2Lj2UJyZC3J+up/5q00GrySp/G7O87Qtrg2OgpTk5/roW13OfTzSvcaDNZ6oST
djr/4wFVoi/BihszZoLbM7mnSjeD5HIWgkzl0ymkofbc832lgqD4dWMKwPzKRrjnjBHc8CNyOHJ/
n1Gt3Fkofk3QqFqB9arWZR+BsmJ5+4Mssjkl7QWwaVcmdIOtoRfWFF9ICBow8SlEKnze31dtbkM0
XnGo4UZ/vXVDM3b7SwML4XUneAYIa8p4D8ErkiSXbqBr9gKy7pBnjdM56ZmK9fltuO5zgqLcRn2M
YY8pE0k324MbtXJg1r8eEQny/CIRXJclCHExj+94xC1VG3skJ4J+n/PqYAVsDJORekJtdpqBXzjj
guMR7IY0ukVZTM05n+GhKSpQifE4InNizj2GR0TqkQcTdyBA8HQPn7LyfsAnYMw8qcDRAF1Zgrj3
EmijjFNliXm8BeF1J8Wnjhjyyx0g7zD9JCSr+ag3W0XfeJg92XqufUMuRf1eqPcPj+Esut/4R46S
PvFcvFz6hnTyK1Aen3yBLuIk9OWj+ZMgJYaKXrawLRxej5r5XZVy6wCEiv4qd0jLHWsgah8Ux9og
NmgKVhWGy21De88X9GC4VOyBQqfEckwmY6NwwoWNKTdQPglz+KuRjKTV4sfSQonLsXjVJLEGyn7j
rUyKoohuifXK5btayupZqPufLh0gVlT476wUYTiZf0VuCzOIwefDvUczCyfjQTYd6hINPBu+qlqj
kf5iHutAtv0J0nCqqbofSM8JfGKVbuKQLK0Gl+W8kMYtpZLXzR3xIO0foWOoRdZGEVvnuUB+Avk6
U3fScYUudWxnze8fq2jNPlKvhCMSOrN7hFyWuNXTSupE5oiFsd6C40qTDJ0foU2kA/sSzzCBr21G
bKwwnnI9ju8IUmHnYWQrVmeHHF5B/RnV70hh7NKNQqAZwBUEXBw6tZkT7EbKIIccKilCiKf2mXCS
9b47fmiqq15Yv1ZJ1x2bvgRAPjnZGCNLcANvfr4yx91OQTWopFTt73uvAmXmzFsc2IVgqm2pre9u
rptl4WAivRA8pPeTdJO+rsyO8x5d/kqqIPDi9r3hvBqASgxVnnGAQb2103NZ4L3PzoNmf4qkiEvD
MoCgu8onkKcI4GVSO6y/8tLXxczweATJCeg//YUuOD06lwkcjm8xX9jMwpjiUQuenJbpIxbqj6cq
t7OfbzTgV+5AEmxSHz/V46M4reKAhdQVSpwCM4rFAO9cVOjxdZEKNlv8p3D97GcUWpR4XnB8Z6f6
HhDVj7zQmGb1DVm4670F1xGs9H2Ycce7458AUW05U/exO5V/25PKswD2vzDXbMR7jDpYcflhLat+
bMdtELsuHmNOA0a//LQoqQ+z/iBuLYAnS+OuMgZBwsjJxdIY/xcHFkLm+o/trGOYixlgHVtrMqfQ
cUESoJIVbXNeOS67B9oHD5fQXu6toEOxyJ5sv+nuRyIc0tr7tylP11Cqa4BX8ISTdqeA2zlCgFeF
ezXz2Lg2CjMhMHDGralbHatgHdGzONobxkou4cpxWNAJaQEJ5jvpUzE7Ct455MBbDswB0+vlpLKQ
BCYkcbankJPzRuy/TxvVQ/9/6yZnLmGt53D6rkClC2UJpavoH60B+ZZSNdyoAosb89Dq1l5h0rd5
k4hoG4YD1rp3J5qS/bfb/6VSpFAX3c5sgH7FBlp7wp5/x5uPKV6mfKW6yqYzfOZpH+siMBrL2CmG
NB1KaO96f9Jq/A7RxZaK+jXKFhNCWnzAiz1ra9HdDvSTeOLxL3J+GcMlMfYtyBJB3ZdWGwKXGRI5
/ncIg0FN/5/8XiP0TMDLDDG2Z1sKJh3RS3QRilTpZaEjWjrVlrvoEf+L8VTVs6FwF5s4Dv8FSSO2
iKCtyZg+bc1Mukfz0FkCchKNIviJlD1+iJRPyqR8YocoT9TYFJkCDs85zGGGdPgG295sCDpAeC7A
gBHDQYs/o+pQC6oNMf1vTKrS1ZCQRkEGe7OOAtiNZJhvQegczjp6iVmcRTn+EIBih8cwtyjvTmXB
TU6zcHExmy2BtdEbJIaBEj4s18gP8V4kl5wRqu2hY2cKAaX3D8B6tVylXhrHaDKU63Yn/oCXefOH
x3AB2nXtn6e1/IQSx73f3w8ZfllRHR6n5MURTksczCCNsSJKY/dL37UN3YT9HRqeRrTy4yLKXArS
UtgYYtMC4nZGwtbkM7Wllt9CYMinyVlhH2L5I/G5S8ZBoclJLLfOBFscP4CBcojcJfh2y4ZBmr/d
/IXKJVNkDuydT01wqQ9M4z8dvI8Fp7xVXbpTaP3soSPghztffjPNyZmpGCaNv1cZV0+apwE/zr9s
kewoMZZtV1hUp95pRUmy0xYuLw3Mfokz62Eh1J/NV7XiX4aIQz4zRtQzcj76Ykq0H9raDwZplC3p
a2EUS1kh0nq5uIK8LRx/Yk8BTVOlqtZxVs7HLbVlGJiHUaHovhNaX9jTnEhJ6NvTVKlsDoopv5Sc
kXSLYWEnzWnEhIM1Q71wAR4TZpLRXv4LN65/x7+DDZOhlB8IwiimzNjyx7jWTttHevtyf11NLlrX
QOmeTNkKO0eUGsN8HahrEUJho47/+Pjn9uKgm3QyHcj2eaVA8+4Tf5169T7v2GXKHVPli5s7e2mM
lCYzRNZRLL1auKVxCphQJ4DFupYUU3bPc6tTJAvHTBrO9Mfi4r48I/oh+QBw86WCpDwGqzv2smJV
/jBmTpeMDjo5fwVE8GCLXdw+oZRBbRfvHrzP4cQJSmoWuNTj6ZRS6qyS7rCuErVSsIxjboxiN81I
0BDzFgxFMHWFvTNUQZ6tXJ/+cbmIT0cQaeVaBlFOEYUI0nyhBqH9mMh5gQeuuxzJaRBXeFzdOa0x
QiGzxz2pLlEsuN6ivlkCSHaWGWUqdnqzv/dT28Wsx90KuXQEFfhXIxceG7ZMJEZXvxYGxWx8ioZD
BDCL4IPTIBfTpavzMLE9PHHx/FRPc2FbTzBk1mILhHroLnq9cnlOHIPCngII6NtSopRcBaa9vuzx
jNyIgU5wUfMWIklxy7bk8SlUcQkjhRShQfyX3YU58lfps4bHkkGPHOHCbnwfQ2pcNZbgT0eXinKE
2BDqIMAMZmH76VOXWisCr+z4or+fNhj8YPfikPadqX6KE/2fMlZpwfZPMLQ/VhLJPuWaLu2Ccekz
qqhXktRIIWSyDlIRgnyLOpS3BC3ob+Q+o4scrxul2FrM7g3nujPWEuMxA9CRDQRl8wz+Ag+ETI3h
riT8zX/CovsIEXCXMwcVjF+++yL2iJLC6l32/FgaLS1rfxMp5xqNlyY4WkdXuERIw7rgSaUzhvh6
vov68u6sisLBHdmqHHzUSL19/qDxZgXaYtcwWT8AEmrYOEdkKpu0jH71dYAp/NKVZqBAgrKy7UAU
T4medHBZ8h9jjMgk8sg9HQMapJdKYSWZeVi55tO99teg63zzyjs6cJiml5JwpsP/+xT2Bdpb3/ln
Fe0YpcgiGmkyREKAoUNf6xDLUMnmIdHKEuyQfaZRtPg/nmmRCiBfdBZcff0l2Fi8Gp1hfHaR2bbz
pNskby1vyIi82Qr4LpdkVJdlnoUX7M//VgKYQFeIA5900Q5yD1vbPYbCSfNNiyl7xpVEmwc5bmyB
E46oIrT443N+SB0nnvfcZGgHgCU/0M2MpaDmsaSIU4rIn8BoHbtIbv8ONmcP1LVBc3Gw+/I+YL31
rXoQjN30Rd3I0eLhCRQfAholyKKE7ZXwsCgaWN8QJUMY8Vj7oQhVx2rP8TK6YjOnwxsO714GCl6H
e9uHN7LB9PO/1dIYIk5j9z/0AaPaILI6gVaQecsgKssie/yDkVbP0R+/INnrQK8n2XkjTxTVwwa0
hSGyLbBF8b90SixmkjKObQ8NySJRa31XAH8q+HeRCkZPbt2e8Xoj8GbyctPH4xs9OB0dtIE+WN86
ihx1XCwcc0U3JM5viwkes/nBNqNxr/PmV6KAPgmOt5n+dwUTOeD7jGTExTpD7MzqCti9zf81AkO8
R2U6YsJE+q7It4pSEeXCEh1zzXfQQfeLTGkx5PnJRLuugqhWeVW6RJ8azZG/bYpABJqaLlE76LIj
bzntuUq4QYWqgOUQ01IYBKZD3tpGgkCgBbltqFix9bMB+T1TYCH23DPtyNkntDuqaYncZ2UAOCDZ
eWGeiWZM+7IcmfUNB1WxBU+dOLItn1S/wEtJGMVPc2JYmelKtq1YlGZjYdVakonyO7PAqH+k6ypM
L/YGEHprrNI8zacYctKWiZpHy+OsjRRYd+fRb56EzrZ59g7N0Uec64jBHMC7VEesPDnsnjFgxqS1
4441g09eFRAjMYZTXjcspsrrlfFUbYFblHVf5otr8c/MTFOX4mev6LECZekKWArl9CF2GBUGH/7Y
7HDGzz3NQABvEs03KxDApe/gKOK2J9jxFZlORK5z5kImbF/RyIQbAQlH/t6PKtNrEUNCY9rS9tHH
Syce88Qz5xJqutr/Z/a2VqxwprzLhTXhvuFqztRd19yCnPkXIYEIzVahrqHdsgNhJtECKGTogEuc
OHgHQgKMQzBAvOvCC7G+lKqWiP7cpXfJevi5OUOBRtKy8V4lf5gRJWBhPspZvhJXlMDVCbMsrEed
37kVsND0bn3aj9Tg5Fc26BzIADYzLUhq0q0mNGCmgdlbTvmqtvtDiXWcfnqoLGag9jZF2rAzYAyQ
3Xkh41GqQe5QD88+Qhf1hXNex20Y8PgsKVdBVuh8I52Au1AYhvHLAkBjwik7UTD3RQZxutxC8cwH
g9/KJyoWFBjyWL/g6lD9l4A6LL2R7VH1bPky7O//Nj2djAJtp4Hqg8RHyuhito5ocdl6uv6DtbL8
s0H2PVjxS33PetGutDtEinav34U/TgSpvoLBtbeOLe7T0DwLmJZ7aKoogm04eWpQVIsFtfByOXvJ
Z3lzSkX/kf7BCm4YvcCq1ugFyJsIfmbwGUkYTlauyPdgC6IimEJfxhW/CXdUQ2R5pf22kVXLvysh
rCY3XjKyR077nLVHqa02fPBtysHFtNwH9wKpdK0+aiPinl+JBGtoEK/rMjFeY+4ptC7MjheR9Nij
7oBKPE53PEWqI0idI4cA642ego32A/xPzf1XgxZbBpxLwsvLMS96Fcb3wxUhNXLYot25ezmJwGZs
7QIYPnPlJnXpphQ1Nvfxjj19dkPaVhCkkdFCfKB/+cIeRiKYDVJG84UVBfB8wQWFQ2B+sXBW/mbX
0GuWjMxmyKW94fyMc51rIA7/7x3Fqsy93McSSQoUP9TuECL4lR50LwL4+L/1HCqzwvvQ9syY2baA
ahmHjfCehoHHZOkKPrwQQkiZE/0Z/eW6ZPo/VNO4LAoHgEdLAUiC8hxh42+2c527+L3FJpbBy2+J
EG6lnt9M9QgRe3wBrpGrJqWYa2xAiImOtFBGtzlz51ohrf9Ss45jREXRwZNAJV82BSiEPJwIG9uC
ePiivJpBl9Gifisia3nx5BwvcRJ+auj6zJkyrSLtkY9cqE8hTbuSd4jfBfSHBuQVXZsUg/q28iJT
XlY77ZzK/TcUBcmIsQEKWPuIxGpNn3oidyjcIpOS2axEN/VM0KJySOeQ4gTnlvmzg8cZeoJGKqfe
rgDYTEVOsjMELsDD44KGPuUYUx4CxfXzyhwt+Hnhw0AvswyvN6iFacjs4k6lWIn/UOibLUWM1+32
qkEFbyz3FBs5enSSSISK/A5rTYNNXeXhhg5vJPJjTSYCdlj5cFCExjN5BIDjKigd9mrNJO6RbSq+
BsrQVNeE/q+o8rNEBI6oR9Komg0hanTzrgDj+3hQ2kI1M5bR9ooKY2T9XvyIHuMKMEvio+SCJTs7
1AZ0kz135aA5FjaLr9BmD1YsTLaLf+82W2Q2fC+hn5G/F2M3IJjOLBFzR5raum1FScdMwv5ErLGs
rxdvG24+jGMtB8O4RaZVieKnwdhH3IIQfMEGpBz5J7/kd0zC/cyFXkxb6ZeLB4kqDdP11sLox2Nl
orrlFiJbAPFiZnZkQLCM2p4pnsLaVUpQRoqqwCx4jyCOAGxQiS2csGHTkWMeFdAMa4U7qtH4wRva
uL24YRzUpejjLfgr+zQgyQ6+l71lies7aGC3peeNo2sYtVPpB1dBK5XTCjX+jcSSwz5/+Rqg6IK8
k1Uo4aLoBi0anuVJy7jl/vllC+eiWENhSYd6xaC2ffyi98IUL+kVPltt7H7CH17acsLKNGhhOLiR
reU/cyh8QW/X/Yk6n8m+ikCVaHXbszFoyOlrruRlmnafsZOZH+MfnNN7FbcB2mx3/5zTa+ULsSUv
aEbz/Uqr++jtl3FzCRUCz793DLy4YPWPRVaSqoC/RkWRXW77L2C35agkLG4QK66BvSXVgVoXvazH
bJseQ0ORzTJ0ihdx8a1Dg46DF365SxFMpKSpXxvYx6oU2mUwT+1D2qtQx1EYwNE/bArh+BUK1zvm
f/lAqJdUL6vHAXmcMFmFmgW7fX5RUb/YyTJijRzeu8hGvkkO2AF/sY0pWs6+gYoxnG2scsM2jTq5
O9c/h2wouWVOfg25EEvsOP18wiovP8QbhzYUBiu9hGrChxpit2nSWDLwX9wVVOBcpSkqE//UyX/l
Db0iMnq1584AXPWeD2TVvAlMSgAQVVunRNSG8Ih3caxff3v6bNaq4kU1b68g7Pb6Irwy3GcyEFr8
ufWLL/rStFvu0Ka5BWYlIIFi8xTs2hFph5jzAFKtZYkik4M6g9Ny8UBU6jwbdBBFJFQ5c8JsfonR
LZafBINYBb+52OXgc7TR+harV4oWmiiTMGG9IlMNGk22IKgl3uxDv3BI31WbzAfcfPskPBSUIRT9
2FwvI9q5gh13YsIEVVXKSR6bycYUdiQnBq60pvb1TNYOHanA5lJnqHY8wN7TVZZpvD7ZOZWUBazb
aaDgfgtcAveXCS1dDE8MNfjgnmu7qZU6YtoxVMj1qVbBgQ8iFmRUmuznBKOIe/eBKs2OL5WGNZOJ
ilouV1TyQaFljkkhRD7La4gdTBneRYp2e3CYwy1wz+lKG9sijPDzNeY1xM+RUfzLPGrFN9uCmuWN
iEZzKIP6ljTuZ3NfycvsXbztOtmWq+1m2E61o8HkmHN2nIl4XjJpKMGWpnIDpxw1tA4zpOL0gmbs
o/8OsQKfGL0B4MPCk8cY8yrwXVWSalSkdQjLcPn0xtTWkhd4Lla/Kp9Ng8J1Td4T+fcIHnvtxqoV
SlmjD1PAfuFn8weO2yawRnaUGd4yjgsZ8HE9GKomdZq2QMb5GzKgqHtaSdphg7KPkN7EIUU3toC3
DIVB8clCGiUbgycwTIiuA6nJEhQtCQZsheBPJCBez33fy2eBWFHSfqBXQdKzTFe1byMAAirAKSve
O0utz7RnM1bxVDhuo14CwuZYalGOpZd1JsAaVdLDmMwQi59iVAMqnF7PNmgbj1y7MRkAzba85BhC
X5WouzZlydIkjeKvccp5yFUYBRy5Na7dPIfV4FzDDUVFs9wGpCqm9OvHs3K6XNDTP6QspmZN1Fmw
aPJ3W07ZzTaFm6peumvOI4Uv8fzIshsti98S9HRb3XVXqVBqkSObV4TgbMxxdLtrYM+ucTF6xeAB
5PQY4FdiOYAqsIc9otzqydvC9UF5LILiCsQTSSan55LHLwC9KsCmYN8QKSGtXT9e5jl3Ke5ZuKWi
mAZFlqwV576BHSJFaG81iAWB24HFOIcEdEFyeALRnrnjjvWQtbWHnOaPpNMWbZuPcmWTKdI0oEqN
BiFPBKehzlgKObjn3Z69ceHcks9Orp4zsNrpk+kyw62Tfmg5zODK+9wy2yBw7SxjrUFcL9tiW2ab
LwtyAXX8f6+5J7iYa3fhRYovY2FYyrZoVLOifyRggEPEqMFzYqeXq9MHZBnooJBt8X9DBkXnaB77
ws2G+qhDHtPYFzlhIPnzXWqyvgZY8iMuRM5phVMEc5c4vds7cEEZw0XIvHhLE/9ErM5RnGOZrOJs
tZq10VvQiWijfF9djs+SMGH7BLY1dsu3iY/hEBwH5qe7Ok2AZbXwVp8xunpdhRLpDPLgzVtQGFk+
+80uZpOqR7zcjv/7Nuy+0I9Fh+Gyt4DN9VJYL/alFzl6cCjCB6fzv4vTslQxd9k9LLZIfYzOx8jp
Wt6zm1mK/sI4EdSleiMTJQEMruOTNBuRhYANlLvFLqR0Lub+e2J2ok9pceoFwvAAlgplHrq1zi+4
SWqIOtTJwd7ZWnORLxM1Gk/+mgoTwpcipJOGlkMUymchmrX0/0FK0ymgJoGWF6L/lSQWFqjWUGNO
SYTpmKYBfFEWn97W8+vtQTkExcx92NUHIN3G/c5y+3hl77LUhGyhRCvFi7zmjKUh2shm/fHiHTgo
uhDk1lpdjPxCYloORIEnQ0XVX2QF19gFu4j9TdkTewX8L2bMquQ0nCL4FKBBQrNJsdTn8VyrbwwD
QnHjqJV0DzU5CNE/pF1LyDhnLKPyoSmVEY63xwaOHJ5gNoq4/C6FYXA28h89Xf3LDAqIj66nELSc
K6eGgDu9lbfVKGb7kGmaofI/EijMRX6Hkt9q6zQVkVHmRoqeKyvR8S01pgbsXc5O4th15nw8Wo0R
lsT0J4B48MLpVuwUCm6Gdb3aUgs+oKN2Us3BCTdaahMQYOpCCLyEzDQpcekkmdSkatwYP+Q8jGiu
DJHgCBOPlORB8i8yY28wjabmD8OaW4f39HMOE750FJjmnOD+4UQ4piMQ9Biqz13fzO30rZtlsYMK
5ZX3LtMSar4nSee9vahBuQiI+XmYmFLRIk3t4GM3e+Ip7txLgwnt99kIa1qmtC2+Ss0n+41e73R9
mepZ9794ZrrntpMVUDedD7EmJci9fgsVGbmmjl7ypjVY6ps4BOg2gAXgpN7lGfCweWsiL7RGWkA2
SXzggTF59/VnSmZ07Y/GBMu6Rn0EnBoG0Xc6kCEsj0DvYkgWWT1QmwI8wcbxO6LobIvos/lJhFAE
UnrR9zG5FB2ZqtUKXtdn669eyG1YX4nXOkNVFfaLyoawoNLJm+I90T4CadKz7rT4uQMfA4KUoLs/
VSfPE1X6DREOw4X3fbiaiImZfm0RY1ilMVeYxg3nueeHAe9GCeg1A+S1NR9kYblprp850asEa3/q
HHPrmhfwPuikyLB8Y4DUarE5EYWD8YjqhoA+gL9fi4w5YMDmg4ODBSMzogRFA5VtLjRe1B/8Q14U
xrmGK3/hpqBtlR+piX1gMfXvKgIBli+U5oQYvZIvloge0Rdx3bDXTxaaD87Qhag1Ow1uzUDlsVVm
Hnu+UimrEbhclVk8Od+YpTEdHpLxexw6n1+lwQk7bpQMIllATf2OjbgufNw4Gf4UX1PrSxZTBan3
DD4tYz7vwcmeYzw/NjDsvzm3Fed6fjh5yj8FAzUZI0HtEY/Zh8sSefc3YgntMciDiqx/HX75qlWE
t1GMBdPT1+0ytUeYPffLxme/1bXXP4+mZWAcm07yiphT8SmZ+xrmUc1GMB/r+0yakLRI7ZP4o5a/
EVu0bsytktywZwvZlY9ZSQZgAZKXFvnHXFnFChfS6kRE3QsP3gcaW4mED7czGy+aLJXysApgIA8v
c/pkFJUtY596LD/l4mskDLd1vv7l0JAiRgFRG3n8tSXP5eoQJlcu7jHSy91cz6vmzeqjJfYzxz+X
kskwZEHZp1CmSzMk+dR2dBIE9LW5e9ARQ3A2Ta9UTl/umXdpnj0qLmsI6/RStZaAjH8pjYXtumT1
kSypqVhgycoMJ2D43Llzcnzvdhv5jL5K1rbhkkgtQCxgc47uCQv3CiCgbzt9aMATVnB3ARzvg8bE
EiM0hQCLeXc2tJXqL2Z/LLoHpk1cbgIz4nEb4CQTicAqPitjLKc++4PyCvt0N4ilXtUcBFqGtyOz
EC3ACsxVAp/bFuvVVXLpEIuL9Kvjx1MijnXtklVN7q/nY3HtjLUuy+fmcSbyV7IoLkkJVJsd+kzX
mjBYe+eXlpsuqe7cKfi3EWIUBR0b524R5yADQiQr4KwzpoMVHQzEGdd1LLvv2h5Fzrs0nC5HMqHd
1a+GnEATpT28uD6AL9wXWA/PumMW3ggxu8I4bM3YpiQcx5mRME9dbS4/TBj98RcfbINsW85DJtXf
Buv3hdzlBFXRhsQBcPo8Pd5wrMflbQ8vGZVV4s0SjQxnRAjT1S2QcVB80uViMfLaQ02IpUmn8ATM
3Qe8WaH+LG+fK4Gy76Q4FT5770uBrpwr5V8VEY4XmBm2Y3vodJFhTG7LPSi6JG/QPkQjYtq9FwGe
phw2AQFMVDeSjHUUfWdguIC0wbNNsFoqzjiszguUXQOuEUocxQq0Kk+Jjgk15GinFxxMmUqLSuuY
YhqXtZl22NGmaBkP+DuTqxJ7QdxSk0qamg+5QDfiODpkl1wFA2XcopHaG4OB3AOCrUlHbHLIU/P6
zNjGaN85nWYDCzci2jiSrFNBPSJzlcOBO0y6UpW/Lc4TADGFZ1kuRFw8vKg60OrHkKbXY+GuAzt0
ciugZ9HZ61kzP0A+eRWHPW+u1zUITLSegHZ330XEcDMsEMrqIKq8zXD9d0N5s+L5yuQTaNWYDFJ4
JM/s31mjFtP7JEoId96rjbFKHb0bMiRMvEuxNr0lgYD5aILznmVSccwzNe6gBiKLzt98Lkiop8Xv
SkWQ/+W7K6PAzgVntz1k3v3ONRu56EG7DY9Hgpjl0M/W9/3vGcKfQbruO3n0bTh9TrWvG50WOaYD
l1T3NDFhZKg9FfCoSze105dnBP1dc8dBICrs2J8ZLwD6kwgtWeijqvLV2g+gXpy0W0UVDdOKjW7P
DI2MU6qHpnqhFqBRYpmxrON+DfBED0vXuVwfkv8IOFTpiCsJW/L4bDlf0gj/wxpYYyH3SyxSN6S3
ZCGlVO8EDlviqJGKMTI0+J16e4Cdbn91OIYF7q6YW79z+2YtT+E41S0Kpf+BJXNixeozw1jzo7c/
F1NSTutXaFs9QCKKRtp01piu9wbHsiPRhWNapJvDJn1A1iwUysPO9njRPtQzD3gRNEqKoy7uSBL6
DyJbb1psCp5mwslZGQAubAWFrM6jnKAhUA2KZK522dm2/waWg5pRNNOtiHO/k91GNtNK/kP2Mw9I
rQr0VXCZj57cFBe8QXG+zgx+LYOM4lBwYizmc4zqM3xphX5NHUhBjHiepEdVX+hCdbBbmT++GstL
0+j4xB6iaR9xMiPy7pyQZ3hf+vdsXMDSX5KYEv2SmR7z/OKEe/28K4GrLdCpO7oPsg6RbPKpwpDn
JJaYC2bG1rByMyOIHounI8HpPceV+6+kOO1NLhYCS1N6Bvtu9JquHEcWbHGkqmVO+Wz9GFycjE6n
HH1g1DunGLk7N8PTwKaMvLTwiXbt2ll6NAByiAQ6YkCphGGvX2exa8p0STQqyAxQsBtQODtjiD90
Wh+rCNdIZwjkO8sbkGBk/wiSqlINO5p1zZ5ocXP89ukR7l7l6PEW4usnAqK1QFCPYzSTc1p+VFPE
OjxMGJcq8ej2jQ4FxuC5Oa8U1AXL4MkX0HQk7dN/jZ+i2b40KKQlNmzBA/VCJ9NuehonJkZVkx3w
pN44zYRJjxnzf/JKEu4uAuvgWbJtbZAolK1/fnAAoinLLjo3f6eU1yFD1A5nU2RQmyQB1kI1NMw2
oOG9Nx5hfkyZYW1+j4JkTImJ4cjwkUj2U1MoKw1dE0PCm1h6C30/U4+TEqpSLJgBbIgGd2m53V1U
yUEURvKPNG/N/nzqhYVRy+fvikBGqWOF3sG/zWK3wptH78iMccbUOSYBMkIk9BuMZZIYRA+bD20a
4iM38tFct4Sii1crlc/ClVRM4oRY4A+abcQGxr9gLdUJiGE4QVyflC1i32v/8+60E0ehEs5ypqcE
2BQZISJ299iDAFEneKAx2xLwipsWSytmZA1JqLjH1D1tD+d1yA84LIRoC9EYkRoAmYLpirgGPvKm
RnmESKQLlccXNIy/yOf04JA8xAl368i8uwRJj+d6IGOW+9jE459OgPOjnFaNKjWeGPsMuYZWFgmS
KLGdHryb9AxPTNX6SBsYOp6A+decaYxfizKuSiZZL1uw5RJxaBSCUosKJv/CYjUWTy7FabBrrqHY
Vh7YfZ5DU7o24v6U/gxqBPqi4oPsNlmnse+Ah4hUWgmuQ1Ci8FMglwa1TfCBvxJZDbAWV4OtpUVE
oMnbibJyZPqKRD6pQGta7dD3Jx11CRFPqqSUGhjItyoBn10xN46rxRvu4EV14gDB14fygZFHnNOH
ZTXjBdCs/wqEAiLSRXueuFyl2xvbyNHnxtWX5zy9fP7Vq6FW5Hm/wCx56JfhnzVu4g3Af+k6Tpim
hnT7nMFeNJMEOX5XxAUTEWnjyvJaX+0K7z6vrMBYPD/sLvSiBEDc5W6wvg1YMYBI6gwkybL60ImG
Nqu8mgG7FjylHBvb2QhoKza5kqQhnpcqURRfYu9Xc8QEzL9rzHAvDqyKLvFQOLDwiplnGb2nZNiP
tX3zFLpdXBmrmMiS4RrMcNrSkMN8g3cToojB8q+EzlVL1o7fVR7imUON8AjcAcawREFLT8MbUC5f
SOa4j3ZAwT684PeWU4/t7qLeE1kt71vBLr2IQWQg6QjRkexuFZ7UJt/NxPheuoev7Q1CSooMgnJg
grQv7//2ApsqatHp/9M5GvuCqAMc82vz3awiVgiun3QTIkWDWYQ+m8DNHBamGYvRdSwGnXtPAF7x
ezuBvq0+arcqRL2kLw5Sb8kKI0dS/Oh+FDuyQBpcZ0smRAGRd/kg3geXm04V3BY+tDk+EPwi4N7b
mD6EqkW4NU6aL6jMUjW3watwd0E/gHL6Ua/WSjTNUg3yeXL6Dh4eBUFe9PZR/dXaystxOzrCbo11
wWCJNLbFFx6QsN0kKaI8AsoAqWaaoPW4WlDbzok88nMhy44ERMIX/qTU8u7YOQ0S2TTIPd0O9e7V
MHBmgxsiuoodvOtI6Uno6BDRaBvpBnAz6vWk9mbHPvHnfIG4XzhQ8KYbbkIVqUpMC2ImMxuPeoT2
WpczjszdnsyxY6sckvKzF5apnszMeDE49x69bCPP5rPDttCFwX2vSnHbp6UVt3Znm1nTVGaeAWCU
zwEOA39z9LCB/wl/pnLQ/4VwtsyvXN8rHewJaDDBClESSJMPkalB8h07rW5IMYGdi7Rqp6zSr7nU
y3/KESuM6KUFFTNk/s2mQxr7dZh7QzouX9IQYWKwCcY8QBfoSuj0xOJP8LkIT7JY+bwcV8PtxKOH
0usw552XWn06EniGo/wEvyEGQNnTC3b0zWh0Gw4RSRNrT3UT84fZwe4wNl965sMp2FKUYSmQLlQL
I+jgNjbKkvOBlDGqYet8yWhqNmiUS/JhipoIQDAko4FJzbK/JJge4UnYYDye5QhU+SE83Q00t/k6
GToldNdJsz6br3LlaJfQ9KjvB+VVxnlOVCXGYgmUe0BaJtEyfuf9jxId0/wT3xLVbkAVDO5ZzMFj
8RQEgIf9w50eaqinrMW81cTrH9MYiBL0J5zmdrTiBsLwlg1fmD0cbx5QH1MdRPdPpy3hiZPJH5Ck
Zsl+z/Y+AhjOkrdqhYNFLqSXn5KYbxZvR1GOqfHxxnlEDn/0ah6j1BxJ/DQ30qKe0uPLOO7N3EnH
3mq8bcp34P80Gyqovw1971LjRm+asDtZ5aLWhkoRHrpn5oqPs0ZWC643CtkbPzVJ95OjpoDmziV3
XraOBf7eQCMfu4YWSCp1g7YN9uPldybag51uqo1UyoXH+0DltrGewdXiWcoZRMVyQJ2bTOKeE1sv
fg51OWFXoepGpjuEMPNZHoHLozZgaPOAkKZPCETVo8uc+grkRp3u7Ew46tdeLzjSfIZGdDNp9mka
rNzeuwn03Y8y4aWnp3Fm9lhZeVjHmcn4KTwAc+dcUm6WJy8T7Jg7Ufz3kqlBB7csiWIWoU7LUYlW
C87B5InrGZyPnMbSfHmA0WMzxxTOhjab8v3neaJP3ouxtSzQ2e7DWxcELAhOvYEyEctTQw+su3Di
CCU1DPX5fM6WNOXlezH0rF/Hg3IcP+QN+ySqxvi8XaLVB7u2JIM4sNFSz7/GK3WS1tsK1DzLh9vv
x9t0WD7zpDFamATy9X03GT4IDbXRE9DW/YPvBOLwiR5sWf23FoijKemGRTfwc7B8frCIIckj54Dh
oJJ2ehcuSprtZaRkapOt5fyfcHqJAKBn+6bTMlF+/LkLwO/PCPWO9s7EK9WhWRRExmUsV/KR07Au
11tj3jBgU7K13+M95i0IfkJSo39eHzBqLhKtO72KWLZsrdmj/8FripL/YbCwFTSdUMTZvsfNn2vJ
cRC6r/eVlYRmdH/LAwrCMnfkWXXXa9aXXeWzV6ehBRd2okxrLC0k82mTwcT0xRRJzOORzJLJ2spi
a06p93rE1cGneUsAmd/p0UmA0pR1T6KoGf2NaKmkaAcLbfyMGolUjDHNuETAd1jxspvUMiGZdX1W
lGqxSO4k1RSa5KG7tOJBzqe6XVAnmwBn0HIkt82yRRD4SBLB9BHeTd97iEGvSCyrM8OzGcBjwtep
rqE0gb3NoEevs8gZg7YDeYurzalZkc5fqt18NNtrJ4L+MnwnwZdgNDG1npl9wA5806k1lIlDiUWF
sftNzI21Oyc39t12E81Jvo8WEkQH3RUjWcmAPLrZcih+fhtodiUhqsO3ZMChFS3rAIg/p3drmmZu
hpRyTjnW5aHAXJUDzpUrRZjSgAg0N4RyHOhrYQzTBKZJBOS8zuCnSPEozxr85P7JBkokgbGvETTz
iA26z35G+fYh02T7sZwffAr+Vzrf+a5Wgq57tJ3IWX0ZMPqgeua6r5hOsHER3YoDy0crbOv5VPHk
P/EbHbVKpqGx8nvulDhkpGHOwcPJa4WDwU0C/McCahvxwovNtFpDKpm3YImvPxSsmqszJF/U2SbI
v+ZUnDGdrAy2DNaTRbhuO3rI5Uw9Y1n+O+RK1G8elOtTMXqC+ugeQkDt9YCBf/NPe4+5PjeQpHzi
aGYO4/naV2xu2i+FKpi0RzbVuZpaIGMbwDhnj1rO6p0EYBWVOCqw3Pv4L8F+o0igMZgXqKkl9u/D
0wKRpNnFyAqK4DvNQauIk+OHrcwYJofr0NPiSwg+vzggqe2WZn0NFmyFDwqZTvUxgmcqAtrE7eL9
3Y7OmlonoVctKj7nr8rhtmVbUVoCrauM4zbzblU5TMhpAeC00f4XCees+9P6UB2865w41jTinPAp
di3kf83V5pXvJiTCePEyBs4jA3A8GSGwZKBB7WcG13GXpIgNJ/Wtl/b4415gNK7SS/MlNxGQ6qUc
IRNujIdf6YBuKWsiDcNTeSunedC88hTGMjeTal8gdEKzjqCuBhpfBHdVJSeZXjz5MxFRHtiRwUyu
v8d3kAZ5lgGS9emzJRzqcBrkSVIYjlbGpscFMf/PfK3Y7jgvZVvt2LHgfFgFi1y4CpMPBjr/FKxQ
k9ebaLvMe5hErtSFQFVbkWd5NMKW/zTlq0vucBl5O2/XlGTR6GPCQaX31BQIH7lv5MuXUB7N8UsD
Sdl2uF7G3yJ90TF91FdkKaCmYtKvpLOOlZk/GODNO3Tvk3eDYxlo/mJ+/5w7hB1gjNHc++KtrQy1
7/dwNUu5OyYsvR8wWgkArBwdhAbm0YTRLsD+sfKlUI+OWNmPm8FY4MN/lmtxIqsr/r2UMCu8wRTk
qn054gEo+OnENBp8MFr9bdvDea9YCA8eugE1mj5yowzby+Tp0GL8zhdIXMh5cJ5+fAV5a408MUJI
zn5UuqWQcRNMf1Jyghr4asMyYErtEBbEDajfUIZN+5sTc1jbTU3NAosPA2oz+Ck0Vu9GFnDFaOBW
UKBEAv5ugDOukC3L1zu0xhTi5EXxBxxNNh9jsondacRT3Sol/6nIl0bEupL/pePEOsInLTsN1UcT
bkL+80DPdQNvuCuwuvvgmVu+0bgr1t061U5pDQ24AZ6NNqfiYR6y+Rbx1kn0vYm68G3f6SVPCATq
vkhWtjymP158L8clrZ4PktN4IS8EDRQzfdG2in80nGCJk+kzrE/Yy02U0VbMB8lw6+Ui/UoDPq4n
S7nZ9LgYhA2S7vaID6qKq7OkFdB3pT51TlYdkulw+VKZ/NzQ996h/OzWGhLO5Cbf4XfozmG3uzRz
hdAy8VrHUkVuODO3yz0UODRaAXg+4NcoWPJ2vYWtNOole9shecIMjaes51EMucpth6xyHThUMYOj
oTHl1M6DNrwSgu0MltZRalWjUk4gzZeuyGTqNqIwZgpZnCwBEtPONmTZL8eCRv5Mbl4oxxODMYNY
smWbn/BiaKtYLRlUMkV/ng0P3948qulgzrasJ8Vd0t/G4HUwS71vmQANprWFunSlGk6ERX3kGP3C
WIDD3gErncSYqgqmFSC49gwt1H960aiHXa7Wp+Q1WnKmVgfdPoAuqCdNM6jA03KdvoEUh5ADVL8G
OfrjamzmroejjPQ70pbRKPLSSEs3QrhYvNKrpPAt3csVTkvv7s5BMQVQwLws6rw76HprcVv9EOZe
zPiQqQET8JctCsy0gwZAJfF8Fdn5o/hN83Ir12y60M72AM6gANUJB05oBcEFurKnQ2zEYrQ7UsOh
5Qs2MZvD24BIzM4QoiXNsL6E0fOtwx4NhE6Ako7iLwlp31sZU/fon9SUpcrxJc/2dtMYEF0nZRY8
qOeripQm1qudc+WetCL9w8CuRjUXVCiYbzENmAxUnE1XNvOJzbXltbsJ00QMh/3sP/PYjwGE7CeB
FiWFav74+je9/aH0+HPbNiOD+73dt1MuMSHsK604gatQwaLbQkxQtwr37g9KygXErhV86Skea+zS
IRxtR59wQJQnfkmpwFrVlOZ+gzCtd0Znr7hTjyPc0wLPZY0/Z7cXP6ye4N9ABQ18H+HP7c9VAgqO
JMqk1f/Kbe0LjEhUsS5jZJuRNH57FzsQ7fFyGbaWe1aZfmXxfgtxLhG8oJcqkMCeEL8/5UlKAQ51
Jr0MGejxMOSLkCEEs72aeAAUvgfpP3ep2JO8zWKowetxoaLZ2PWOo2StEnrVr6CwTda7d21LWahs
GfaV6PpDh4CAXB8uFjMG5JuORLQkT9XaAbnYVtCMzN8R48d82RvL4QXlkPRMqCPIdPv0GFwdsUy5
q3a8PqlxerYRnFTvZhI9rIOAvNkWoObLS0/Y/cxPohnokb7a/ZQM2FwCkyrME9roecgZIfm7PaRq
RConNFxGht4fBjujSFVf/RPg5Jqw1HRZDFpEbXk6GJWI30k+lqWWMsT4HUghi4NIWs0752+xI9VI
D3ERiTvQHOSGvmpSECAZW2i6SIza2jFscDvVpyJJ2ohBtbR+kf6XOmRT5vTV5kb49IVpan7AWm/a
Lc1upolhsDhw7DRdLhwj4bqq1QrOkmkx/dEbptWDBIsNFXnJJGzizVOiEQnizyDlsr2iOAeJ8irP
8itV8OGuAtnwujxzY35NJIqJTQGWeqJLaiys8Mw7mVKkmmNEZDQOtRMmngHNFwVsj4LAXk7a0s0J
FFwm5OsSglEWvyhKQ1b28thuX0L67R5XNkdLgRmO6TqZ5IO2dtUZRnYGkXGUwlXE1KvF+rEb/ShP
9uX9mV7QYR7dH3xSWvfKsmy1E/ReS+bjnohciqRxmdYX38vyGdyAE6UfAZR9Po2sHgxEzVocwrTZ
C7ZWDhO9Gq1N/t/OxVA2UybTK/z8VnK994NDM2BeopRYmyu0P3GWrOQDOaCs0lDMer+vEVYVCtzS
38yuicPyEmuhggda6h93h0T3RQpIx69RmjOsfOaBnm0gdh/IBFtRX27JQBNcpWdLko287rOl+jwW
ORkk3+vwk+tvywac6YBqq7mJzZWj7lGkkehVUHaJYERIXT7evsb31/XKvpxj3kcV1whsbLokGTyh
Qh5v3OkiPfA83hJY6SuXk071oGS1fGXTwXmEJUpxxte5eHMbnbyTTdEGkmLI77zW1deH6uSOy0+l
w0BpymTCTluqM9BurI/VoSgtRt1zD1Dv3uZ3JtROoLgBrgbdMd0fW6ZVi2SDbtmxtzTgAAqRat52
IbYg6iKW0BDh+SE82EOEQu1ztSpDhXjzrMPEjqFVdDdTr2xjA5yBn1x7gmHNbnVpTItKPpUtXk3r
KVlpfMX3kBrVcdlQ03QtcsXnRwtRLM2lVsm1IP1bCTGRNi8cxoWTwO3F421vt+lfehMohxo6Lm0T
RLLG69snk+GTIxvABaNvaJ+DlRUaShIX3/M+XK2Wsu8lFTx8qWOMjlSZ4h7onndOcY8q82GEHSQR
EwRw+TVhrNrwsbIH98fZHcI7neLd+p2D+6m5imMlfJgS2mwxp75psFEA8y9Qxo1t5f1FfW93iT5T
nQkf0jYaz1+PUizoJw1w4Rt8s8LpQUp1cJEekBkCS+fHUidKKoyr+NG1V+QpHosi0mF45pnVrkg9
c0nWLH8Is2zri6yUDWigGR5pLGPT38pdauptYdk1RHL86SriIBvPOMs96IF5a7ygJ1HDGjXC0cby
De6IVZs9tvmm2GK0SpHumaXAvtnj+PFyk1yKKnACXUlcO9iOq2GSoV5pd2/Yh6ItLKbE34j1yuVy
RiAJZhK7o0juI/p9N9j5Ax25e2Nh4DSsk0dooCA9Xb6fC3vDPjWA0IyAslorI/nTuj7W4sMPCOJE
5ErMPwvscQxIzaSlVEE1g4nYZjUreFFwaZOZJrB6qrIqBSHKa9bgSDA2SXS2NyznPqrADdn7kdHu
gnyAY9IZgYbjJwUyya/ssOw5Icv4ckzahppFZGxYwc5DYdYYv2hbiqHKK0+NMcQLaxiAErSfZ9MJ
/X8vhO2x3i+cQ5Nv0mcSMW1bcpoPALvTv7B/4Y/o0qQQSf5atByseoZWpmRG9N9DBSp3ukXbc+Vo
mdoKSY5RUncY0Y5enwBGiYGQFRCtDygbkrKI17zynSZLjIKSlpqG0FkTku1LafBlj0GNMgYLa0+a
Bt/aeUwNf93sV9tm92UXuh0X+I1ZW7JW+IUHrSqLjYWEZ110jTIwEGO4XxGjUQtZjNW2MJds3Inc
9pHL1G8ZokivNDVMKnna4ClF4LdeCBlfnUVw7aQTWTVvi2bea31Wr1aF0eSDSskFOciI9a4+sX9W
Zub14eSenKMVl3kO9UDoUKPTIO4+97Y4e/9u32CYKpBLC+qNKJICbPXq0eVa4nLmtAv1+WtX4mWK
pim6tb6XDKAtkM0X2y2N+MV7n/jLUiJvHDbxzja+f25n+HugMNJ9a1U8/KynLrCwZwJ8PT+T3ycX
3fkuQdrFkoXPDW1LXh0/EFB4Gz6Jzc+HOir5Wrv3HsbFYMsZZXFfKfE+bTd1JMZFJQuGVyqUqBZc
JfAJ6fGJ3VBZseBKmDe+HKH9ThAfIZvWo/PN+hq9p+XfmA2pP+BqZFslDgdVX9z/Jj9ww3GBnSRC
pc59A5lqPZBzIvFZqb0POw63dQCejGKZaHrmtLFClNhxqudWkL3GKxoTk/zMXEgSJShZ215kJkTa
n6pV4P67nL5qMVA16vgl2GhbAYXkLqv9MFh1aJ3ElI2JduvkYx3b/vHJvNILWdlMO2FR8fxJW3kH
fcFcrLVGJiX8QVoLbFXGkaLTxM2W58KXsaIJknXvhmw03+UHUasFVGGsp1hdQ6HU5RXIRRUX3DRz
x6fm0vLlPu5XIyzU/ZB3dDM1HK1eIDHat8fNGvq44b8gRnfgbsPAEwxp+B+UNj2AW6IX0E3Nr4GX
4flIO45Kg/RNc4+dvrmYgQcUZ3QYKHM40xoiW73wzyrkzWNlt+STfE4/m00C1YTc9SoctLbB+J5M
FVpBIxLwbj6E2W+GSpezIFFrwRkY1HEvJDRJqWp4D4FzlS0FNI9H8aUtahlLCXns2PvjqhmyEThU
B9IcwYhNQblwgHgxz190bvazOMDhMViZahTSZckwGwVqWHsr6DxkxlvOHDNHBqoeggBxV3r2929T
qk8d8K7geQ+XXJElFw7zkgvvEFuW96HifPKs0EmK0yDacxg+pms9KmiWbDx7PfsVy8XdhUAcaUwv
CyHs8rgdpZNjBUCMvpTYhP273mocN+hlwJB5jZJGr/r8UcBURZy6Lr+LvhrcOczo6kef3iy7TkdQ
gJTp3+pHIvGCjbM6Km0G+1v5ULOoD9ol5OUHDS29u0Y52d/6azYx4cUK9QVRyVFg/nZzKDeCXRx/
YczsVcja05FJ5O7bDHXzPW7DovMtJW2Hwq/HO8wWXipHk2L1XaNnsZ6TAd/82k+QXktchG5zKaoF
Oeknbiv1EBy/mRmssCQUTH4m+oHUP6sxs4By5SmqM9Qgq6Spz2i9J3TilxZRDzDxvj/d1gnBBGex
06P/K/3iv0gC8EYojwb/eyGh5tFdlyDPS84q1Id9nEgw54ltSfD4g6pY/GW1H3wl/OMVxZZ1t365
My588zxlE4zm4yKUCKssnhfvTbtZwr8kl4/Ppv9i0qTtVlTMKkKatXyXcuQn+dUTTuguTrLnFPfp
XZzXr4A3nGTxTIFPZvCpAGAF9EthtiIGinV4QArdRNSH5ManwY1bENg4o2IV3DoEkMwCCjOLMy7A
Ih1lxU5D5PV7Ms7BYUFNkWWKjpoXUpPJc83DBOK4oN9jNg7wRCRM5ckR77mWSGOeA+p0URkOH7qt
GHLGD9C2CofLVGOYl37f+iuS5YjyCrSAyVnrBY5k/xrKVqvwvHHcOGXe6ZwNXxzATYa3FGvkd4UD
HFh9k1r/u2BAblsyZGrGgBcAmoLyamis+6k8YC4KMt6W9oAhc9SFDsg0BfDDDSs4BYjO82+SLqRL
YHn6R7JpEddFGogMRTJt0IUrCFGDj02jqOIRGce1KOtq0G+oFXndstDIqwCrKlm7Byn9htsHY2GN
uiJGn8Vj/vyEUCbqKtYjjwLFS7JlOvjSg+r/u6EAbgHaCw0SFbsXkb6Bdfi04S0J9O71bi9Pkci5
OVYPNWYswcB92Z5+bt/6dzmCcFppPrP6Gh5A/+DhIeBOEAE2UKu9WEc3dcmkeJoPLGNYrzCSjlH5
3SieN2JKLsIeQpkR9DWShJ5NBNdNl95izUjaxlH1ANoP6gZs6QSiyFCYCfmeR/aJE9CqIMh98tE3
XgN5qzpKh1jm9qJAEEd0sFp6REsxs86/z88SvOjFE3bB5ETPJ88rst/agq052UcAhSdSvDFYWF3B
NJU9z6b+tEqzzyf5v3PUG24sAoMBIC0ULVgZxT0PtwVhBrmXv4IH3fD+q5QyCIq9kKOoVU96nNXH
ecI6BB12vu8qE84a94YDxPgNFh9iy2I0Pz5+RDds5vD/qbp6TRZeTcaQuF5OYdNgP4dksXofiTE/
AqTMzg9O9aUlky3CJmauoFLXl2Go7gXaV+25l3STUKq8xZIgW26BH6YhhU/Fzy/0DzqcNHnNNKdx
gHyA0skN+dEnnkXBKnG06XHoJha/uNLni1rJbEBtOZMW5JYIKl7Qw8ZBob739F1dQEtQguhMrhLm
EE7wzfMcxZcbhlxH9uhrjiOfPoNPK+4oKqDUmV1jDg76DXHsleoK3SgPQ1RWqda++ppPaZcs0SXG
teq2rDKp0e0P1KYoLKJ453y16m2hXZPOS+FuBqcIx54Jlldsx95W1E1F1Ges0auTKrhB3R1HV982
Gj1oBPtwysL+vZyJ5cEnAgi6r+gDUUZQcais5QrwwwrVKGZpSqF1itECqZKMT8jqsMko7M70EtcZ
I5qOLGwcCDhLEaty7SXqnwPvNa6Z02yGHA0eriYR3605WwK4XY4ZugKtau8A4IPrkFeYNNNr2eHQ
ZwYIyPA/4wtbASd0oj0bUk3+S33ZHANTEspKD66k6ux0e1ryhq8Ta5TAFHnUfg8Rko+rD5NPO8lV
dFAm6JhTcgB8kDdUVFyv0OMMacv6KlL5jRup0ZGEggUwXWK2YBub1tBbB+wk8ndc9kD5kEsPQAEn
6jA/SFlfOxjpXivYY96GU2psrSSiWvP8CYvNreLcKleCCMDgnYsvVo+/ztenY4HCWb0shKdUuu8w
0bQxspLukTkRXShGuvqxG3nvvEFP1TOOTlI3qB9aF5OnA2uZkYidieY0vE+Aogep1/GHzZVak/0b
rMxKnnsB56ET9CCgme00UiGj4bdp/tU05bJVuju5ipFcodVSMsNaXjxF5uKddCVnSeU0aHZHGeH5
U7hQaoK7gXJZMYdfJ1C7VZUAjnhrEwnzMXlbPJaZTUg/SEmlQME5+/MJ6XJZbgfv+qQFlunPeEzk
M7vwVN5n9MR/MlmMdIwW35QrfnKBdo8xMQ7/rsx9Vd/RlsWs6s8l77v39CerU/STWKHTpEP4etfP
8gHes87IB63I/ueCMJ0A3n55T5zEyr/MH7O4UR4PgeW4nQKipNc1qWfaWn9/+3YVyvRJMVpml5M6
2ARt3pZ1RBkiHvQOi37isKqHeNUB7q0rr/80qR19HIFcYaGCNYSdHY0LCW9MOuwt8heX0X5CHjTQ
mVln5lJmM6/AHdOrLM7YJ5fKZSj26lb32bNBNwjVTnRTgoTjLZhedzhdwxI6VDcAgflYMXmtb93F
S80vqmpLfGI9mH/fjrKw4xmyaeFS3wIPhKpxNBpSAQ80tLMhzLviysqF3DG3ijvcK2nK3t4M0ALl
QevEYSrCZAkRv3Po9NFMY7qcPvI1+9crmS5As81gg/W/6EaDosOWQb68+peOmeHoFsryKw8R/Dui
TkcmiFPEYFZTwj+vWvQgGjg4VeW/U3bmCf4LAp7pNQBlJmXClCvPZc/nW9TWH1spTaYo/PzLLpqx
0KvQBwVghsHbWN+mnba4mda7R8BRpxGAIDkxDF2o3htofEPWu4VLfs0EOr82KnZdJdoiMHH/MDnV
4QkN0Bzo8sZT+q7j1I4m1wd9IO+/Emcda5120qZNW2Q+dBzTG3fk1r9MwAEVFaMZlSmoOMyzxNvA
PTEPPraBSEo7KAJWe0KVwZRTlucJ1UDnYhUTSOT3CZYAf5JT4qne4ZY7DqP+ZFlEkPNr6DIiqTAZ
fwr4k3V0qiPnpa6xHIYgQ3qtwTFQEBl2/ek7+EUNZz5nO4GqQxbgujwUa1BfPH0m3A/lVvnzlMoI
jXS0V0B/Ui5EC+WQdAEE6XaFmXZIJ0PzQDHpgTnZA3Omisr4xG1b6TsrfybjeDaprg8IKTckd1Xo
EHDeJKXrDvMlWwTFKVff4FLBzbprrHt1xWymGiyo2mfUVnND4yl7xcmYagBobfr09KRZONfr1Apf
WX7G81z0wZzSR0z4kZnvthBQHV2qq2dtveTNDT/IYEXYMq55uQ2uUC+A6ddk0SEkG569QfJ1gVqf
8n8pfUdA7u7bV9jkL8SK1A8sW+GWU3uUB2oUUGA1crTkjCHH4pkp2iJUDMEyY13L4/tLQIqz00KW
r8ahYNChjZt7afKJo34h5pov/83BovB2YlnCq4hApnx55erucFufgEgpR0NUJH4eBMnXaRcPXFpm
PGeiIg3S+cnyPp0Bi5uI1UAz/FI7899zXht0PEptmO5Uhy52wFyjHzsD9thJl4R1m1kcZi1/3Cib
pxme7DSYqjxjm2eGRvPs1jwB3njxgAgRSw5TsMOcq/TFaAcLkYW3ex2HMKX7n17T+A6ExnNXFSBN
26wvT71jL9PoA7hTCJ50gQpMz0eFkS2wdjpa0s83yT/Mz2Vw8UBPpY50BVWpo3ckqrCa1vVimDiH
UAtz6afEGxmFvKOChP6N8P/LKZ7SoY3KimXRgNp6fmqiJj8drXjbic4OwalBPqAvoaiDUuQRCnrS
iMRMhpfqpaLRUr+/7Y9CM5Favad/wRdA6GP2f85Xh8jgx9R60+PSZlXX8GfDKe+5wHDHLpNEHLLd
gczE7wTEOtmwZslySGfUYCMtq/YU73mAtX3AKN6J8TVAAwZwwiGtUgrwzTeIqpzF9pIr/ZznB5Ce
z302imyL8YxWYAGcozBudyIoXW3mm8HPU9wKgInX10rFVBJm2uhHunzcEHq2ZavQo+kKjkIXRXKN
jFRH0kOHqadv2pBB8UuomgRqQxPDYMfi5ESdmG4bKqCY+hvgT5y8w7ubTCfztAaANi8dlTtVDZim
Z3otb6isW+uFuzNH77/fBPzWQ16GXzTds71vqHF9Oxv/qs1fcL6VhzdGDVqIxFGCtX27MTs1DKv9
6HiCH6muuhKBI/uGTi+VFmHxs4rmbG3lAwuzpq0BnP5cz8Uebp0QRE8t9D1uns0ow2bD23OtuI+M
N4XE7lIqgTX8XiuAQp4BVdoUpwzoOQdDiac85NKpmYEK2FiAtof+6ha5QkgL3GsMvGSr500hNf+t
eZjN5sHjYvIdmtcjiUIVfWUJpZE6iL6Yssjb6w+/6vxUrZO9l/0Sx7LBPY+C8GGRR4xywfV9P3f4
Pc5J1VdxrYDYLNcwYJYOkkncfk5DGe4QABHMYEOyA1vDUxl9AhuG0EhzwSjTCcUhH8oaOj0Hzfsg
BTt9D0YvX2JX3moWT7gjvhIfHK3+Fb8iCpifnUvWXuwJ6TDzZavNILi2cuV+/zliGn2QvvYDWj+7
QuY9lL6vkUntPRMLJH64a7cyoqwtNpq/7VbddNEEvsE8W3ppb4pInUHy0EMQi80vnh4nL5px3GdZ
re1JlCIm7Bxr3L+07t+SlIzocG+E6GBXEt9qFPCph4KPLPCQLkh5ZSRi14qv4ce5/O7iL9EsvU78
foOtpn4YaF1hobDPBwcEIBQNabhod6gThgFtdAMmGRQEaGi9y4B7WbQBKWNEycJ4uNEsKDGJeQaD
Jy+VHK6RMxIBAFxYvJlatXe0BJVSNOeozbIbUbuzO8Zj4edSDIcEudV710j85QjZG5je6ouWc1sA
1dtAgg+9TF60HkVgFzSoL3OtqcuJeauLPIa7X6stdE5iZeBLP0p6Y5tkL+YZ3FC90rTFUshYzlmo
ug0abw80lG0PrXiWts99fKecLKoBfu3bfD9V06oImbDqMj9CSlRWakKNNrmil3DZQ0MlvvW4PSkY
AYJ93GuoGrSbwrP98OmMyWQG88PTYx7fQhop+4nFZrANcrwPOV8BALbCiiRYRlqhozx0+MY/zVRD
CFLM3lhjPJH7pLPmPBmIftmUMs0QmRjfXxXtziJCaB5W1TS4+CoMsL6y7GIb3OQcki7kH+kgj1iz
lfJcb39lM+hKqHXPNN11df7e+H8D/XwDdGEcq1x/bLnUzCyxF16vtJheV7g6uBA49Eumg/4jIT6i
OYdNkqCztwcZSMkJPW9xnazBpqtmavZ1yPVRtsA/89OJMZqC3yqL8Mlg3Q/utIpNJ++cWWfqbbi3
NseIeT9wMlf3mflNZ+28BBhf6AlBnSNmW5UvSjWEoxVNaWzKRfFa6uj0J+gcK7xeNl9N8VEHIhgs
QEWWrbu6JaypoO+LMKxo3YewnJyLYr+O8pI9ajl/K0JPS4l0OKBEGqgkWpPeJSZuzhP1W/14IK1A
lwU2d7VQO/5KKgJjIkuBaCupKCOZc2m33dqLpC+IdxEeHDRJoPq6hD6ZnwplrHlIn7M4peCpbvAo
GLhcRK+Nw5fH8cYjo0iiez6VgqXpe55ARYcwemrYwzMxLaJCO2LcIzhSiawrEYi0pf0Z6ix8hrNV
XxZol0XNQPrwDPTJtTt9slJvkNPWCuXchUsqeAIb8jFfFoln/kqaeb+AJA2aANjF++BSy4+Z6e9t
AG7E/Jaa3ZEHVrW19BOgEkn30eTBNXIipaxmALr4+EEDG/1w/cnXw4ADLNEcBJE9oPL2LOtYuPDl
MuDPUACHoYSuPcw/geqd5RBCVR0vaupNUjMrOJd3ZkOkFBbn7y9oCcmm1ty4vgb7P696+1QDnxuk
UX5bMqcNBiJTHvQkXUdqJ283PmL9iUyuTidvcTbwd6QB+iFegUnipuyx0Kufml4MbUASLNpzOVQf
EpXDkTcWYrtc+w3/Fbe5GZrptIots2I86eQy/2gONF/DpaQ5JTozVxFDPjRUZMZx5HudRTq8m/GU
QPJ4LoF0kyXjr3P6SLgWof+79WbXRu5ZKxBp/DdtMB2OI5E1RwFhRGZiz6EYMoATRH2TDBM9BV60
rfsRSpNhxkIheVVrR2imgg9pM5EhXbAna8hiVPXFwoOeX2JHpVADii4eFSHqK68bH/29DAwdrppp
/AErWBvnySKBT4vRQA06w5SZnTsZzgppvBbL4O4iZM2PxxBmd1nb9zv1MMBl+HvscIq8bSrLODM7
upSg//POjqh4pHdaYHkfDcv++BPIADElcMX3xLtOfpqXIf2+qfzLcRdQxcY3G5skLrHavXMbjPK4
opCgagXua8v9eNT9mvjPJkGp5nsJjN+E4Ky3DUBMcrcdd93Mo5PvPXwWPKo0CH7MyRmcQ2jmjjrK
e7qXOZLFAdF17YKNoj3SYcesKEbz9iarxOzoxov1v9OY8opDXpYbd+vTQ5vm8S8ACUDCKOA7iLdr
Npywp6qlrhmIDsb7G6hHQd7nsPauFyNB9JWrmQYa0G0tXryyrFHZZOLloxtaxovXVLx3oESEGmjF
Ps2yEeF9ios8aW/EyRKE8DFeCzOj0XI2Q1VQ0txTWh4GexzGFRauDqguBBFT6aPL6dZ8Gm3qSLIC
sHJ1FFIq3F59ZBS0SF933Dst1QP9m4siKVjDl1ofkqqvGivuCdQuTBkAXudkJPSYlNIdak/ykTk8
dPfV0mUX+FxQsRnLKKyhHP14ZcttmHiclUeAZvdNhg2aig8SrmeRWLuK1Mp1w6t31Zolxk+JYdsU
xf+l38vF9HepIOg+IghYPox8xsOeLFOliD0uctYebWQqD8+YiWoDyfzc6I758BEv0ABIggRUpIaF
oCVF/R6uIcbFmR7IFi267v/POcxGpi1ixxwfhk59aNFRNIjjKRLVnb5HWeJz4U98kkilrfZzsgwj
PPa1hYI4yTUEPu1X39+9msydjR4HUsA4LNB7X+eZlYaM9FbSZYGISFm1IpG+2EXkBXct4pwTych9
Dpntjcht14yRXAAmaE/5mH8d0hyScF9SYbxEJHpAF+sTisVp77jGuTXwPWO2POUrnEQxIUFRwNUA
kmo8o002suQYB0TRL7LFVRMXaLmIGerQa9zp3X2K3x5gMtnHgFNe59n3o+/PPh5CyCGbShKxN27u
23vR574oUDptbCaX9P+1lcU7S+0a22OCQB4H/niFfJzcz/JBH/tbhqDJPc9jQJ+ydWa/ZqgxX7X8
to8rJ8P+ynRb5ZuRVPl/sdnI5TLvVmSsyBJmamK+KOdUAWh9yaUmjH1oMfZcYsBIBumY7DI4yR8L
U4xQe9yN6m5YUQDex3ewmvHsDZMVOU9Ww/X153zz1aijoPgZivA4BK2uU8yQFHNEH3vqL1q8kULr
EnkxCTTvhCiGxYBnzgmFb2kGQYfypkTZ41MKAjSMBFoavnzz8xRvGnbcqTijk6U3y9TiVIzPGcfh
8IdQvxIpgqxe0faCGFNT0qoazDA74a366y8xk37pXM7ncDQKqkOKK+9bIE2ae4L9b3pd6K9Y5A3r
435DL+l9tZI0O8ATvJ0mMzqX8BGPGJpfKyfBmAzSZiNFADLE/XF3vGNJWwQvrPVCRfTyrCQlGCY4
3WQNClnpVcIZidCYp2RQ3p+Dd/lVEdIAxfYJSKfHi9+MZNoKlZovif6X2MiZeLksIlBPzEU1g4Jf
2j4VwJdZEMqQ7BmqlHeamEwQqRyCIWXOHu8gUQN1IebbQyzIuvWxkyfm6XUb2TmMI8jFVPoxPHjk
QV1eJI4C7uzRZ0vZcg+5r252FBnWL/rRtsIkzpHpPCm/UbBSvE2fy3SsrWsy5ACPwFKOrZlJBYLs
DfV2wRRVR7D/UDcWoatQJkoy2ixD2KYXvDSK/pVHm/MTkHDN+IZtAg1SzVO9Tm6YTHCGfCumUw9e
1YWkevgGLpsDm5f3UnFP7jzrL0EAkaFB7pUDcPi9ND3Z5V/tNALI3lYsVBQnbQJszHFryCeJp61d
6dmMIxSUg1dnkWv9MR/69MFeGUBCyzOAsEnGw9hrRS/yZluM97W1iGlNVSR19HyTXuuLvmA0TvyO
yKJMAwiIfYF4CVXgewEZBGq/qN6LvEFILx+pPCE9ZoUby6D3O0cFXTis662jyEDzE2AUU7/PBKhG
BQCQkxCVeQYjjd2/7M9qJJuN4RpTxB7JH9NKCoIY95kt8hsFULiDhfpe7d6DlpM8Q4twA4I/8vD+
c7Yl3TIDwFVNZ0sZ4k5EkaTap7th0rfyjpUkODlV8RhRIKlg7VN8L8NH2ywDyOpVb+fuvkoPYKfH
meF/oerlGkFS1Pl5upzrcFGEF5H15PfzBSCh9CKBjaNtAgssqOjyf7zghxrSA1bigjTmLYbebA6r
Gd+hYq+xRyOQcikzQ4KOZ8nZm4pFTo+T96xr0GOTuCmd5Oc/Vups+capzhb1E8MUv6CSt7CX/CNZ
KGnarQqQgpw3M9XBdWrYmN7AClPWEGmm2VC//FDcN3sSxSfrLV3Ua6nK5rCUSl3dpTyYr0MQPTN2
Tfmn+MehIs+cB9kN0oPQAZLIuiUp+9S8Xf6PxE686fbRpMV0O9/L1RTtjs4lvilL21IUyzVFrhSa
CAh9igzj+oDBRG1DVOWReONGzxulfZWKcVtRuEYHR/JgT58OcCcavgz8eQnJoe0KvoXBFZGTyUYp
Y18XmsitsLmOZQfYQZeD4kUudiTvYZ/xf2iRo55Rfyzca+ptM/TAbXCrL/1CIIqs3gEOctRhcXTx
OsQs5iNwKnWXN+KYbrAYjrG0fwYjhljbVdwTGQW6hU6J6+xrEj/y7Jigl59lDwKhpLO6WACfRFLt
1FFFckvuOjcAhehT+eRg6sMVj4FcpjBoWN/LyjQtWQ4N3iHgQD8zEHuS8pXKRD8nulSXYe1Qrozr
7ZgQM8XhTZARo9NKtMiV2aMRwEuFqPui/mugCQ/hDC+NgnWD6ZXOTPVcijeE/ITL/ot0saFGMJZ8
t/Kj6r6F9xgtovO6oWhXAZ9Gv0v7rvlFYr2cGboyfVJVyR2cJ+4ZGm0ePOdX7EAeYHonv/iMPsPL
5q/JczUX15anBw4nphxYmyvJFRXE7s3MvTki5C7ETXM922xWGja7l23vBQisvFM5a1VEheUR3bKu
JPig8GqUWC0ub/9e6yrUltm4yokmpKddVQSRj6XuY3jvpGAnw1v5j5XrS7YWZl7Mp3T6X/o7c7e+
q+lUUXJIHnYyLCBQIK8qsPcofKfTzgVIiyoYmgZRC51ehlgcLeqaKpJiK52ICYNYg/ZyFVAe32OA
RDqUxCXVt/71aYOlQVSPsWP9JG22ecF4Qb5DuWJIE9cJ99Q9qRw+4MeNKhPq29b2nLF5bG7iFMvF
YbJW8+CWxuhcqGpLC6YtU7d3RdcJoJ4vUIYVykAEXKUFjGDEISuiWEYEwBeZDPbxHH/8vDNS4qP6
mYSMlk3VQ+nhvlq0i5qutTNm1UGxi1VjO2M0O/noLwZp3NgOJcWAFZ+F04DifOHw+drImLVVHBiJ
TNxb5NMl9i0eZWAfGQLqBA1iGKfjQiO3cqpX/AUuT3zFa6OOlmTkY3jdBJe50A0LfklIdj6LQeEM
c5w0DpXYUVJ1lUx/SNcgzf648s6KlNHRsNweVS4caTQ5DHr6QwvEseb4B6JKT4iUsm8rfJu4XmuB
Jv6rEPreAdSr0tNYgf2jucH68jCBgSC0VQiWSx0njfyY5yiZcbPxQn39ME/8/toP9rdlfs+6jMWj
DnpNz3bfxnB1gD8Lz1GxkwR3iFtH4RYr21WPQe9ENfDB71g3dBUqEQnQAsoj0OJKP9IggfwhME+J
vhiCw4So3ZDyzxQmTDArRtX04hH2BUWQEV+ckYkm13d/uJRXQ1JPeg/PClhR2mV9nYLL5dcKDxwZ
DJpMJx+oXLKwHiZp4+1Vks6SKd7IhTH0GYhPTl9swO+yTZVFzw8P80MMi5jYHWPQW9QDQ6rRPRoH
Io+cDboJgB+TRIxY2hrDz8uijSRYQtpmqZNXO6Tlo3x8de5NwUqK2k0d720QlD/76TfAUqeO+E4O
Wj9UvwYEv2pwXNF49N2LuX+12vZigOk9/8QyWTHYtwbENCxiQhClY8XqIw/oXHbrrw17MGpluEgw
USRKFH5wZTdmP5Pm9Wj9bEhUoD6hoYI5ueouy+4yakxiFTqZanZaVVHy8w3xHfxRbRMoo7Lxyxp5
0YMMkqPMvFR8Cq1Gxud69+CoV3CnRQw92aBadPyWPQN0YymsnHzjVE9NpdNswjkRSmhgksIOT0Na
gyxYay2A+fBbDmnCEi+mVzjvqRobfk26OB5o4+nf5Hp1bgnJqXYQ2U+XLQi+xHhEMbkQEPEHKkBq
9U3YkUiyebs98V5ISvMoLlemZURheyv2E1IDG0ibzm4toOrDN42R9oWq/WBwt/2nXID4BN2jUC2C
hUeo+oMUcAwCVR6DMBgwFq99y5wd0LeO4v8GVOj2SIJvFGQ1+1dDeGrlfYwxVKoBpLSvVCFrNH4h
XvRRwPKolm6JaSZvunx4tizoHnPLIUupkJc8+zkajnCU5svoa5G0rVcBn2cSU3gWXm34FzQhz3gx
NS8c/KZc64Acca9V8DkbXuaIANpNg1o3koV2+wOOpGYbMBYF1TRuRoHiEfIzEmLV1XUjVd77SioO
JamAzajduoxgVUHMI+NA2bK+N3AlahhkoiUoTbzZtmrlTQ2Wzf96dOIiRREtvA8fyfLMuASiijq6
oCuQmj+d88anecH3fOwdkkWkVSdxbN8JgLq+mxy8NbL2oHgP0zcnxycSWC8VmOm4hWHrCiVe0nt6
d+hCQ0IQOAw1aiDgNvKYuiL2qyPL3CrK5Iaem4z15a+uuQ498yAgWlxcY2QJW/2F/MOveRhVO4qG
Ee+A3ZITtmfIXxIcYZmCi+dYG9z/Bn92ohylESgLYlKkyOS2De7QxfSIPR/zZA7rYpiU+EMs513Q
hVQjTOIvo2PFH9JXEXZDBAcVCUmz42eHlzB53JNWF02W2dfvgZ9QjGR6UJprg/br74fmLhJVxfa7
MKjY0xz7W7GY8OSZqDIN98tyfDLNpY0B2KAy9ocLltHe80H0MdDFIC/B/HRk2jAnLgRdTG/cMwGa
9rATEtyTK3Upgy5wuw4NTLwo4xi+p0d/tWosdt8xDqFJ9wyRepcmI5YeGs6Vq/NdhsjwDiKSD0ob
yrXUNVIC9vqjw64ZNLP0h/PF7hN34y7OB+UFyyF89Z31oQpNc78FC5XUpqsDkuDoZLoMLROMVBiw
zLk1T2oBIZCKahZMz87hT+hoxgSOoHheRpc6gwj0uJB+Yp2Wu8u6HOvfYBGHmub5EmnUc4Ie2RCC
+VYMHchbwQSvPn8twwm/DM1DQTXeS+I8f+XANJqIlheCjmEgRcxfOl/4J6FJTlNspPFsUHTkld/3
cQ6dEJSMTwK31ir4M68/FaJ/BFqGFL0UpNcVbgkdglv5oAwlHh/fUb7iSAFRE3furCjF5R/Kymjt
vbC/M4Df3apmVgZK2ZHUxy6b0SGCnY9zWVu0/amMSV0LQvcMo07JsEU7aM4Q2sYDQAeu9KSBjAUN
rx0LQdz/M9p5ZWatM9l5wRaaiwU4b85cvrl0e5kXoL0ZZ6PjE62vnlwXKVU/30f56OExrfj6bhRx
eayLCXDzvoSWKcnVNca9kIdE0kHIw0Po75VIvVkvxhph7HWe5XVZV3pISAqQdfo0jEea6OyCJLKi
ixNtiW0kGvbiGvep1W7Rj/ztwd2wPP4nuxtuYmm4b9MmQFlQi7uBsirEfaZmmZ0ZXgFE7/rPOD0e
Lg0RbisElbnAPb0GTyHDPhDzq1u6U2y1I3nVSo4UNAPYtycKErhgdkvwIAMMDo7spY2+SgHHi5PL
rHY5AcIFm6pjz8zCpbkghOvq8G2F9ssGv3Adi0ZKCkp5i39NETZ5TYrZIN3MK5TWGfSuplQwKsbN
cjfTMs+f/VGudq6pUeSYtETsW9stJoD85npq1H8TD7y/MPWiNy9R2iNsWiRjP0xBws3qSTdkWriM
k1ZavigpsgdW7kiPf+N8FtFiuiEISFN52CJdu8T42P5Xg680E7FEn5CwP+WXrOlcdUy+8CiUE6Tu
XcmX8+SmA0izbQc1oe5hrGMLzwVf2ntuP36rfrVoTDt3dV1qaMLJPRjJAHird+GcuPcUFTqZZVtp
9Py7KoVKTz/4uDlosRGvVcAXHnbK/xF74tbQrTr4DhPBdWCI8Lxok/NEy5xH3kQczmX0WUJbu0+G
oMrSJer9I8AizKyEvnnzFN8urgQFptkN/CtIH2nFCWG9dqQj3EW6K8VV0ygi8tzwxRmO8fveGwQS
w5vfkmaLBfqVQ/RrbEtb9biazd0xxXnkCyMhFftv1WNJrFvo1Bk95kDsjpmuaKpoh9Jkd8Ui59Ed
Y0g9AJcl8G9ImpxqVWFjFG/jmXtk35YXVXgvU4hqYeuTaPyZqNh6iiYb1gCNSkVR9xp+RWKRY7Zu
AnOf8//h8gsCXWzQFpHnSVFsFObnRgh2Cm+M32kVY/2A4CKx9epbtRVjypS1E+RsEouNpwP4uTvC
GBZ70su0wR7svr5iNlQNI/v3LS81oWtKIxbIuHOMeegR5ep42KUiCusLy2PUElYGDILmne/APIPi
YcCUViGahue2/8W7t+PAOnTyA3MtjphJ6wLUSTNytZ41Lw60b5G5zFSgdNqZ4Az9KseoYHRfJlCW
0e/keZLqqb26vgoTMoOJ71gUWsI3Lo2S1gihXpnPMSohI3mxipjAfQXD9WmKGACiDaC5oGQ22MS2
4VYQSqqCelHZI29ccLNzXzGuvq1uMs34S2ZWwVVVbSjAaH3dvl0YGOBzDgx3k2bvo8Xnr0vFhB/F
QTWGzc5JHiSypmCPqqVok2AdNyjobuzPEynvAUQ7wXgkUYiD6BdJfbOEBScbAViLHWdAcBLLHfSW
tAfnvIRJwuyaiR1IvozGReC/yiPIyYQ8lXlOw20f56n9VSmRgZ9ZzmWGIBxC5JTLyr+kwUB78zJG
WSn20pOK3HruFhosbFYcKjT4H1QHQxh58ZgrLoalsEK5RnjuRM9YN6GUS0TnkBZXB5c0JlNVwxdx
LwdVJsyFpDDl5OR6B1ep1zLtNJ8+b1oLZoy3vLvg1+V8PCoO4NCJHF+OlqnILUSda55k87h6kop6
unfM68vZxKnGaa2UADAUjF+23j8IaMPpFKjfDQ1e+r4iDJ/Pe261XnKKdFYOBkvEFvUvOg7t1hFI
CYzS56hDv3UFnO9ohl87oypbcIT6+ynxTBaym8KyORxjDkZ1Ymz5u3ZVoKhGkeqX65QOjzX222l4
Uxl+7HKM4fYHbKExmI7Kcgmbysl4o84LN3RrHoTSjuHXLPwU6Jnnq1I4ry09wn+HdLNfsOrI8m3B
0Omt6Dpmocrh7CigWtnTLSRn7qOfJ4Q8YELG8BnIgBl+218UqWYujsODVaNmprEGn5sw6+qIfhfg
OAQ9xTVI9daK7DsRvmY8BODi34zgynTg5SY3mQ25ILy61oYOhOAA5QnwM/BiRDe4abFrnYKQnQxZ
T273YlieTiRqZcg22V36zbj+Bsh3vhDPKTxbhumaGiPXbyWxiZlMnmJ0RlCfyFO4GbmtGtKmPUeU
7L4WzO084WM6Ex7EGoOZyUlrONfoAiMqtNG1I9Xx7gl/r6tsCjXwlyK64D/kE4o7+Q7ruSTVfopt
UGHpOZJ/dnDYuPBI7Z7+u+I83tHVvmAt3N4tpEzngl5uxOXjq+CdsHXhJI3W5Zg95EIofRqMmXxP
1QPYtllK4h7UeUpG7855w+4piEb/Jox7Ja57j/WFrKy7UjmJQ1H04jDb5PhuvwJz2i1nfyZcY9td
rj7nE/zphkFzfgsZN+wARK9fJdQA9083a/fxqRbiPjGaGkECfJxHz0w69eOIlj41H/HJ5PprSx5w
9LcIaDc52vDM/WUOIzubvpIes2l8QujgkU1aamY9Q2iLEnRluaGOzOvC/UWoAPEouLwws32jimfI
WGPasdBOCwiziIk/h42qd6iYerdNnD0x9IKjRhs0pj6GrvSPsx5XFcqFJCOsLly7R47tt+ZrB4XF
s59IRsK7BeiCM9h8FJAgyK93fuxigL2SdxvFrqLvEAkesCagbycATu5MBVzBA188PnSr2rkWaEFQ
KbaLKpLDLUiDdGn5knBfgvLJWp8LeZofLnV/swIuPZQncIGyD0hTZraJGpBNRn3DaXwBooMxZeLs
pihH2E5xINaANMzN3heTy8AJVsTSBnntUr4Y2sAMIRJjlJ9D8YctdtoTILY9ev21aeWFlzVORXVZ
gpdszvOotHzq97WtpS4nZD3Y8ZIfFKkccrHaoCEAhGqqqbzn5HUajVY2RTaOBcA8ozHo0K5wvR8D
cTkW6WfwZdS3mtbtCgqh3QOYqLsE0EL0a8ubTEJK2qaDRA3J376MYLAtGA+KjPBZxF2/qupwScCh
5I5AMYTyVqVEn8/nw2nJMz9SwelfGmVWpZtVzix9jMPknthmLoOu7g0qQS7a0HPttAVbOA610o8M
1OHj4DQg3Lwy2H0eUY98DTj/tOi3WJi3/r2EajeROf1PPP5uPSnkxP+f7rn+6vHnu8JFXbCCOqaA
EaA7pYJuLSZ12UNlAQ1StvDbR2f+SCASNdamkazMPli3hyFhfzSo9buKo9abGBynSmp3kx9ZKi4P
5uTVQv/6voUVvM2EdSXGKV2WRCG7qeCpHzuIY/cxVwAo2ZRnbREnzXIKB/jFSYqb6gFPi02tuccD
ZCU7qWGR37oGF+mD1TTs4cj+qzpCE/xf70aITz2yjLr0IROCm6NxrBIia0X67Uexzupt8IpDHII8
HGzHFR1fKDXtUi77zNuSysN/ffjaQTN/NK0YOpjFqBQy+VguFy2MyPn1i0X3JpEpOjd4sCjjuuIa
JsIGaOfOz+u/cSTg8CU/NZybA46fG+DkneI7+JerCi4dAijNYB9UW4KxB6nI6ELJttvBSEiiEeJX
E+WUoW/8G9LlLcagVXIl3bkaAYLu66/DpYc7vRqgb/rsQ203APFsCtRDm01LDEA4lxggksc6JEB7
rCjDYUcyTkcz45gpCvXhvfP6tpKCCSrAWLhuVSZ/ZjLy/EKqtZ4jCVAyKyjCnDgi9cKG8t5Lvamg
89hr+HEBlsmevXPXqQQdGHtMKTjNf72sDvu0zaXv3CTrProQOE1yNT5IbPi8Q78KNgjURhGc0UGJ
fBIXUP+4QbMwi5Qm8mDoxClpWK8LbX5DVNKdpKcGqP2lo74P2nV9aoykls8K/laYVxlXpJHt47xT
G7mcKC3hsCVreAQRMTjJgWZGNMBc1LueH4o51iw2aTWpbKrKI7JZxVi1MMb/XWmSxiLAF8bEAHWb
5bDAMRKtFtlo5g1MgfDT+g6f0gRrGvckJGpabnF1rPV7VlpeffKdhd/Dgse0VAC2mvwd3igFZibz
etqHGkOXPd13u0JI3GEIXBPWcf8tishYlKudew3ltEE3WSVFJ2GPEpagKvs3I/h00cy5dK0ecYe7
idfy6ciwQMGeuvoUS9ByXpYHGY6WgVho4Q7B0byW8UlI5gTOIEIiD/Z5onbuQKvtwQ5bUMP9UvTo
x5p4W/Pnbb6/2KtVsIdD+IMyUwijnMXRoH5Ay2Qm+5qi9CxTZNEmgW5X01znvLydCkUmg6ToZElL
HFuzcYbn+0UO+TkogdFm3S3cDJatMrGoK9bkKEcpwG1JkZZrQc+CE3NY1gjZpARzrcAeuoG0XHny
ROT1MQ27Cryb1zSbRot9Pv3Z+DhLRZ+aqZUkaC8TkbZpxJNtmhA9AccII3AkLIyti7dg7MZn9T9g
F0xxKvwTESg89P1aSl7oQpBTppIuJKks+OA/pkxYdjhxsJ6AGeWiljlST2VgS1fCwtAbzc5RxQoJ
P2QHyB2YemwOHuZdLTv8/Jn8f6XPITxoCL0ZulZSCARV6sIqoC45qKhFk3kbcHflB/VpSMGqva7G
Nc/VIQ9fsM5+HI1Khu/FWaII2XKo4BGBfMdF4j1kdzgiSw9Uv+ehisa+VqOe2E/T9IF7oItKTJ6y
vXmNKyPsTGOOpb96o3Yfw9KES6kEe5smDZqJ7LOsGqxQWR/W8da0JYrxW/8Gq8yIEx9TLLHoo0nj
PpghisaTb+e7CszVTHBABvQWQC8gduNG3UVdF2MDRDkQMnHprBk8f41I77SQWaIWlikZoYIbrgeP
CvdajQWTGiGuWshVUOiv4R5ysCG+EO1TIQ7qbUJkwhp2XZtPBfyWn8vAJcZ1rSqXzxAr8mHoECPt
5SJMYPx5+FEzIXb83vxhQH+SSOt1wRBEo5KaXc1A8lsFS/uHR8YfHNVmavkQCWrKJPNIc4jloNkV
u2E69T1CgviIFDfg+TSCoLkpKRW+lHudPDTrSglLUc6TkTp96yj16NX4CnmpxTcr9oDANeYhW1Ab
ZptcxVciKhQL7k8LDKIp/7LTYZiRT7JScQG00GeM4XXMlEbcQSfnYbQcjfv0QGRCGoi3NlEFJGhS
92AK5jZXJuCdDBjfXyPHqgblUJAfND4bz8AV4vgf1XGaG2nPYUd5u8xvH9kBqG2+JoqTvQcv/s2I
F8di6qtjnjF7evfV6k70ajMLzH2lMlXdDSaTT5Kz4+1pxxv/2WqjFyllwMhMSJHbFhkOT3uRIsaF
Y8KpDrWCIl7mPsxcvk5LQgDd02Krc8BR6aCeEVXnVz1dOAfSdcz/0tPfaoOERRtAaY4FbrDpeCLk
SZ39Yky2Hm6zcFmrr3bimmADwVVvmPMvAY68/6Q8kjejWxG1KqvoeKA9y0vcUhQOpMeRkWl05n/R
krMNxB9hTGijV2cEFDCvqtVjuyaoFxAycJigf8QALMy1lrajwSf2DKxzoB2bXIcXrbr/ZQttuHjX
cCd6JY2wo1LDWtLvlly5ABFwZft8xeDyxNT2XnVFtaxxJrvYK2bo4GXGOfvNOgABYt6x1EOzUp2u
77C5wTXS91wPSZrxbxt7v9LiJqnm219D8y5Lk8QoLlwJVJYSrAGM60qxIBns6Nf06sR0sGXvYjT/
AeVcIvh4WCqSs3qwiNVrqj9bkGQpQVOjamucHNHMblR2tM0y5dn98GUW94OFHR9Hz3rIvejAxkDW
3bJCkB5uzH3MiZqc//KdkcoQLysfHFaUu2iLd9nCa5olvU9c7BNYQu9z185ipVqrknsvK0oD2G8w
VijpmRZl42R1sTLKSaOYsSXJefooZT7pFAVkIA6fH4ynAJiQYrNXEVGSMNgf8z8EIfKn80MwsCxN
oj+ljy4P3mrqoBOiglv9YDZX3WQSKKnaQ1otJQHUSH9M+UCysyebvE5QTmTNKMAsuAh+ad8C2KRb
PtBEKv/nUVB6ol9oTuyGc7vZYrION587NVw26ZKp0en5QMc8THEePzXW1fKbHcMmxb/l2gLgmGQw
G8aFp9T06HuZn3MlFafPy+Pw9K20ofYAxsrLfz5CZcfx9LnLdqorawDL89GA2su9izH2xxSF9yOL
ljFHs1ynRFiY2y+LZ5/oHKGHEmQtFs5dqyeuqL4av+G/Ujxh8MZQQUsjkaYahXmH0TIo7uRnlCke
pjRWXrK2oziQe/GfY2kGcrBwueFS1iG6XqcuxNSupgO+j9GHlQEJfgZAoRcdwWADWbxWwjbfuLgf
GA7QnD/igInfBTJI3aUnNbEe4U+SPPcVWgTir3jOsyfeonyWwYObi0/IbO5JRaudhVYWZ15qiUf9
Im8kD8w1WTQKEyZ/NfDC7VsEYXQaoSLEeSVsxzqQ1EvbTl9lydj8UKUGMOG0NHmjgBpR7QOXwM0P
ILcmsH0PtoUyASYLiONTJOsrsMfPjsxi+04dd0wwMn4Y2lNgC5yuK/+Nmw6hSNGMvrWMKurrWw/f
l4PtHcovwNpP5FxKR8nBdrOsGJ6nxRv7jnZeoSHarMDLEnJ9auWyPNw1jPEjQDKQA4/No7TXsCVi
r8JEzzmq46SgfhwFoTBLnIOV7G3kGJpir3IevI5iyXDxY0Rvm3d4+gkk/CJqNB7Z8Ri9C85eR3+/
LAVrNrbWSE2yWaS72tUwa4JZXMRbk+W0TrmIpp1BJksHSyz8U3pd5T12IodXhrKj2Lo9688oune6
S0W5nXYmOQbZxTtagUCRCD24jEyLwbyG4KoZJemfej+LqVhEsx3PhY1zjPdgHHeknhdjRfBjvhL9
FYDn33TLlp9danGSgtHh7t7BgjU5WCReL4TdzvtgTMmUPa3qzZy5Psw2uPA9dc1Sb4QwT90SHaII
ldfLAQaYwXhcK2Zg/s2BEwDN91P0tyjHy4dB1RVWMG0rfFJpTeBeeelcKktYAccgoD1D0CWkdFL8
6uWiZdXx+YucsErlvlOOf7MWrDNA/TDqNiKqvEtRTrBe/xMiXjDsRA51IoM1caHiK+82+nIWDZ6T
He+wU4aURkKiM8AYCAqtx5g71zCIp8DZ1stW14Qrr4T1vUIDDBrciEc9Uxbv1PpzecwgRMjyNxCU
bRu9vv5gAXlxlox/VYHRCsS0Yw67QSlq9Yc/jPZGkO0OI8ssSuF9EPcylS2WZecHJXU2RpUdtg1x
dSEuuKBhjeWMf81+dAN/cEHvPM5NKxN5OyCeBAXfUTSfhT980M83NfcGgiFe7nNVQuhvlUh58CRA
1adiQZ1yMscuKLfD1pgxf4r9IZu5Swmts8ikvXkze99wrxT4FAgMYLKAclKgo1FOmsQ6A3DOAAJJ
sinyXz2GLTroIHSgb764dyjITeADl0tWVvL+YGvJrdeYWoFgCg9kxQnnAezSo8dDFj9QpZPEtqxJ
sD9HJ1/F0wvQe5cZwGeds8j+UpljD6Qm7td9Kmq724tez1V0CUHwMtL/8oT5V8JKGMd0EQS67dfl
/bor/KFjmtc6aMPPfLPa9CViroHfPtRtud6xypogqJo9dsfV6priuVVogJol1Wb1agBBH2T0RClq
3JOxuYm4BH1EsbpF4rgFwBa9xJSkVlheT110OB6OMK8qOYyricbKjPAgX6uz32bRlTCTO8+9Q4LL
hDfpBMlBZq5GtoQIsmUq//+0og3gBdXq/cMoglkjI2nbTvnhhu69q2IkG95Hr0zIdh+jdv/4Fky1
6i9tr/hJ6NTmmgy1vHEJDK1d/x1gehqRRQY6TuKGog9vjBaBCC+glgz3czZEB7HJhJwDn21qdN1W
e41AVURKnsFpgsH/aG6qyfQF6m45ZHpa+tY+JqjNhfRg8iLoVWTNyprHzKsaFPDBPuA7kl/ja2J0
1pSwkgaVBLmM4x8K/p4J8fJ4xQAFtuxgRrU5Sm/tsrbCLI4IhjBo8IM3jahOeY48J25N3OKJb4L6
Zc1T95XqijI94yRXNor7UsmZZrYlnVzizlqEIG0Zckrs/NXZyXrywhlMcSkmyvL9hJ8i80JaW9NL
pmjM7QzQq16b/kISNyuM88BKkhyPVLCU60qHLRxN/Za6RWuSJF/I6SEVg6jaz6GfqY/coRLs4lY7
fNSUY+YQhwj9dbAp3/TB8sVYfqkTr0AWEG4S9/HtsLlTnzEVUp3bbKC/TFcnUPHJHqEA9Z9+wc1+
+cKpKYG3f3/xeSScfC6PKA8E3mJTtMOYR2fYbYmUP8yfclzvuATgVl0isMYjicbE4fU5k2CmYm4M
iouscDEo4Yp7Sa11PpYlwA7ciBM3df/7kLyi6ySJj5JCwBosVng5oWEGr3heVsgImTp1uWP6AzjX
xzwVzAkWKNBsssZqby2SbhaWq0m3Dapad1zvbS+s3E4YzhR3mroAX9lnmRkf2b9oqymkUH1Gcz5d
nv1pMvQrrYoXhw+FB6STRaEG+i7ThwD99HxYqzRRMOKrsW5mrizxoK1JR0lTDw42OtnuQTHbRJuf
MBRFs9aCph83gkFE3HIrw8MCouHooVQxyIukTpjXOrirOOC2/1zzTK6in+Fa3dwH6Ekk7GM4FjDU
NTabwTxIMX/siw6sUjcKYs1VlQOTtdeyVZGMTMMjreiWtGdQm0TPhN+sulWFPUiFUGlrmxV+W0pv
4J6p5TPErtf6dGi+Z9TjvmMC3dZ7RTx/Lb6psjZMWhafrvzAYt3wyfLJVSKisoJ9fpnw+8fyXYpx
tUz9KXX2jvHhb8g3SUB1h0QA8RV634hdcaw8u+nL96yHbdcjgXeSdcQo5Ua4Y30OLH3oSxT2ttWL
2VDE93MUArXACfMZWT7GGsRYUiKzorSAJ5axCbMtiKaEDQehIPRpdz3Hq4na8C+mmciIxYthxUZs
M4NPn88cMnjIm0PLNWp5+218IhZEED6fLXCEfPaasyIOS90SbKWByhynigoJN4iplf1zMvfLjcmC
jPQfw4mxYXW4BQBb6zKz3tWh+2LnKJyVR/wfrkFB8MDG+gm36hBqmSekCCM50bs2aN+p+vDO/Nse
3c14tcHRMChaLZ75+u4XaxA72sJGHWjUcfQrTHRXVc4CRvAk1914owmWGY76vmBHaemsYrbXquhi
SzdROFtzpaejtKFLc6KULuDwQqJeGUSMAYd7ve5AZnlbHpIWanffAbcMLnlk1Qf7geMOoakPiWlS
jaP6R8ZZnIaqfF6FQ64iPqcmQm+dlVwxJ6RXFuh+/dCoAwzAYjkfbRPTv1SDpX3c/EOLRZ09fv0Y
KrxAz6li3RqhwxpeDiDGrVHY2tOqgBEhbCN1Ci5gCGi7mPLuArYlyAmyjR+UZRJJrmBdFdWvTlKM
jm+LRvLq8+dOykQjxyO3o9RHNRMAWpy6e2TqUXhU8uCPtMRv5pIYG5iutRAG6QYFfFXfud5VXlur
P9K6/F2NrySJYydGhZhGVR6TYb8/4oyk8N7uU2h8GbPqsbnztX7d73ASFe2rqOP0qnXItdd36+AJ
zz6+/t1bEqqfIdNE8MjTesTsD1k0LssZJEheS+eTaBTDxeQqvMtKj7LA7YU0ma+k8qNKRXWQ5roN
ojcFyWj4LiawdVSu2rmzSAdHItHmpTj3Vh3prLxt5xLp3P7ml9cEPbkllV0R9DoASnBOwlGFAr2x
PNTeNEj0Yo99WEWF0McTZawPPiwmUPG1x1IOGBbKzd+BRWtoaQuhNsXKUQk9+iouN+X3ENZ92cff
f8EbQyTlLnKYJR3txE3HrwYqUz9gDVxb+uGEZOuCFu2Lz5iKFcQE0hw6fSsG92OWyb2mPSvk547W
2bkrMwOP/prf8Nb8chwwAqArKFf0iLd/PlFOOroIEU9yMAksFf7W0MQb1IgkhQJ/r6BJcEZK/3Du
eadxHMRTbtZ1haEeeuK8/rj50dbdiFKB+uTNNWKfL0/2un6rKcmpfJxE77QpIE+7Iu4ri/L0jOoD
Nt+CLuDch9Rde+FywAw8zf9JPLzGQ+n+Nvrq4ua4qcWtAANvl0q9bvyJ4sPid7mq//PWiOsYRFoW
0FK0MllKrvqdID9SMr1nfFszNe6687Ln+pjYPPYLk0AAranS5spKvV4OXh+j7HGuM2OW8Vubn43f
HxLnTbMfi1OucTB44SpkSSlWJQzLCuKJKvYRUNIiCHdLeuawqPBC749O3DJ0TVnTlIhRpH8nw8J3
mi+K9h9y/DTAjFpueiBCPOg4RjilBr2KQJWwRZBPS1uMI9zxHK6kG71KH9cMUEZBRCfqZk8K5wCn
l2noOq+OUAVQEzs4Z54n1aRpfYOQCKnESnGa5cG9dqDNHotp0wwcphGqaJgon3ZbvAmggh2KxMCQ
PMnKvq9ivvZFVWTmrIWkAwufJ3o/VurRSqzxrZRiyaiQ+trsooA4DuhX1E+ZjFjhEH+Q69ZfpUoH
T24ukXAVUIVmb3QnLNicNy8U32xTEsVzEqlTuxBeB/36l2ztwVaImk0m6lR9lZeveKBkZhSSYiMG
blDLUpuZGXUxqblH1Fnaq8hCMsDb3uryQG8j6crd+2sNk9p8FuWxV1xQYaAMNdWm/yDhBUQbpQNu
eMZbEFh8IYLy4+XNL2c3FyprbVmwaZKoZ6ylM6RYbCpQ1ZziFhxd288tkcseausuHIBo552KvCGR
N6d+V4nMIpaaCvSFhxrIlK9TWsCzYWRq/7EsPN1xYB1tlDpRqPUb8mnRroAyT9QBUFAsC6eHWEvi
NVfnStJW7vLei08uXzKYl5536I06Zn78L2qkUNRCgGpM1CqsJVcvj1/vCLkJrBxtVcE9+F0hVUhu
eqRNUnZyDHA04oyXb3lbjJGgX5FD46HkaARhmF0f3Vy5U14iJEMvBpFMKtOE4C1vLAqHv6PwOViY
jeZj3Yla+rY346MGkHqlAWC4ki578/v/0ql6XcfIwJ28V4GH4MlSMwgdzdqBAnhdEjiBPfwxUdEA
sAws4cdkWC38czIHH7ard7udtfIyYtNHwMpxtAADV3ImJmLkDhqvEzcFtn9/oVMNQSj//WufFXWw
IX34qfi58fdNv97a0lp3zHjzlJd1P10PU1l8DcgeneIVln/VgSOVDbIu0L3A4gkyP8fuXyVWABWc
NVAmp1cgcysHv25wWSWatE05A49PFglYBR7tDJEPJ8zsK0OstEYIOu8MJNFVMX/DgigODrCzRijN
Z/TQgVdLMEUveVRyH5HYy7BjflAaozaLnyvGOEJlOYAQN3JqTbkSMQPrbo4IWPPwv4jdLP3VxHHW
qcH8m+/G/BzOVaJ4+eJKBEgxglOViuKH71OjE/NwKZVM56Qif3p5FaqZns5iOYr7F3JZ3kekIq28
DNaLEYbpbcY18gusLeaUz8mOgt/e1kI6TieHkY7Yzl3DYfYkIjtpB29qPf/tjG4An738VcnBPRye
jrh9i3UQX3h4xOhe8pqqQxnx1QIX5fKmxdVrrXIsmhJt5mHuedI2HxezyNz+CLT2DlHm1fRJR3GM
dhgBSrxXCyVocZOjhPdXJ2j50JGP7Yi1q/AT3zdAUnSA+G8JH34BCC8LPwu3HZSx7C17T7dQSd0A
aZAWcfl76R/2mrSitlPMYaQj7JcfIhKhmV1HqTA32IVmVesmUyGBvj5adEAxemyJuJDrrlVKTnNa
EPUMcPBWhWIRtCvj7sQjKtrlZ/Np3lG2TG0523EFPPlRP1RNa/z+0eCPPO8T/mQP0VMAYK5jAcSD
0pOwUrQYq6FYcX+grUfUo2OPQkJ3RQHPIFO6X4cghTs67a8zWTas4ELYiYhmoNgDnMeietkiVThH
vufzvpKuK6Oe+eDyhSIj9oycufTHh4Z72cvxb3wM/Q77YE2k/SsuxWciVj2CbVqAV0dyDuv6Pbou
OLOdn4ZN5O0+IrmAzR9tebRlabgXnU0ZYX8hnudAm0C3SaoJDsMugbdR7D23RhQzUxkij7Fhdz9W
eNBmvsdXAHwxvY8JaeIRYeEtZhVEVl+yeUPLr6J/vFaG88Hq801r54KfMP8sBn70fP4y9+yuVgOI
0BMGLmtcRb7s8Hxlr4POXQE/EsgcbFt5yDCvOZ0G6D9iLzInAympyMdZPJNhZuzfh52PxRGOHQP7
qOKH+66XGbbXLkOGOThsnoOQKEaqF5j9OQWvqwOMwzLfXqFwO+yXz6toXHxasIM284ukej9ic0xH
bHirrSBhS9ksb5UCzq5aWkDx9D0lW6RaSqkjwKmG5YggIbfajgP86l1d8LYQ/RZ65kfgZGI0xVPC
PhMqRRuHub5F9yQTYAAlkZkD0dPd1XlTi7t9Dl+cNY6zhHIbOP8dDpHefCOqsniV8/aWcx8dtPht
4mWHhdtNJt0j88jWg2CME+X2KGMySUzCi+0hoUP+i4QEJOVzZmkW13270LcaOGzM8xe+w8fGf4Dm
PHuRZt1WYW6Nxnl8989mF00e09R3ex7eJxlbnye4Theev7oyM6717RVl7aXHX+IywPVQUNvbe2nT
jjYzL2GH/8GRstOu6S0ZpWnVqirnwA+0M/UXdiZN4n/PIaNgRimBZ4RF7xeVYDbEjY2wer+ZmmTm
hifqSI569PjXzrv6YEWMnE+Zz/ufAYn8kG21obW1CKjRz/Q/6FRdU+D8dlVbEQcJdk10zjMzHwaT
b17iSDufP6wzAdHpkvFGo1aI5qYbz2NgsPt1J6KBZ/TxReU2WWt7RS0DJGeXRAWVpXkIgJOimP7s
7jGmoht+igr3V4ECjACdOmdsXik3xU6JRIM+32l9XmRnrwo2H3udtjd2BzWkkJKbzSnshxbuIIGu
ADK9ThIWjOLZzSjEkHqQYzsX7IjoD1h28g9SVZnv5HMcurNoVKsgc3JTaF6DwU9/Fyx7h5B+m5q3
yh5tUtVG6oS5cYQEfwA6EzqFRyWHQDKCCwogOI3tibkIxEYOGeTBHFq+5do0teUj8Y0rffYbnzfe
pK9tUH4L55XpBh2xXv/ZX1N/0uHMvQI8qix6QimXXxCz4iAiBQbUKNCQoaSb/Hj+IRdLkqhA9Fda
YwTTO6tDZ5yGNm7x4E6mHcJiXYqLw6MZZUBTN+AJ93p37o25/I/uZiglPMPzl9YU3HkLpEUcLlqj
WxrxVIJGXcLbl+wRqObIU9LvEW3l/wpRy6hQTJZPYC/3driA3/JLtvop71/8KwuqSEVzOGlDt76k
FlbIboMozCgP0HPNwECjiiMGfIIRt2FHJJVlA9mGxom95GOV42uWJ/MmouYXxvRi4AOe3FXydpQS
zJwkkijqLYA9VkdL1fjIx4BTmt5Kp847PtrcgqQC88tPlJ/Ty2R/MJ36kEJURClZkrHnx1VOp9Pn
IA0z/kuhWz7lsjDUwie6bNkOiOcu3scmYe1F11DZHt3f+M7iX9eGliaQhNN73WYndZ0aum1Yh/bp
KJQYnE8JcOmF53wDMHSfBsCdlLtbY/naS5TIftEJnOS8F5Ez0agx+JwYpoYIPdIjmp20Xx3CwLf1
BLPVILJbxUnnvjHy2Dv9xpxqbAyC5adDFp8KMCcIYnQxurMqDxlD7GIQqi6rdNAz+n1zTe7EAJMv
oR66F3/8Xv8a9c67YuFjZDr/Tmg+/d1JKPKvcSQKLSSwebrKumPbpf5YL9zfShKBUC0/X1sCybeq
WkqiWcGCDmGkwnmC7/6eVAW/7lYQHOqViJXuVGLYU03v+xoeqEO5NzkgMxv/kzDpmsXScLNCzRA9
G2nQVoOclSqujkVGrME0UD1cOozBAvUZCCTFU+HsqwTUP0U0aCiz86sI5S3pT4s4g6POMic+BWhi
pnpuf0xe+johruO3F3lb/VzouTq51mhxzvgqmAgKuXKgQnbwttl8gbsOGDYSRipnnbhYb2FGTlK8
F4AdQNNadghiOW1bzf2zZi65KMbOq+3N3CSXcbkrICrhELXY9u+2kceF5qLYae4QkjWyVQngpu0k
4O5mjiNV69ioxanvUhUFr6HbY+5muLy7Ud9ZlaQPCJSWwaueaKTkk9mq54pif5JgDYvOeUuVXHTV
tNneGEhJixqZAEYAvLe/2mGnLojoprbhSRW1dpSM6u0Q/NWuY5VWE5cajhOfvPDA+5Jp55n3a1Wg
x2Yl0Du5PST1c36g1H2jMW9jmtVk1OdZNGp/3RCtk+hPhuVljEQ0FHMd5RFh18BgI5wr2ADdZpcO
Zq7aSAWgRLnffIRlblf9f/x/Ihj5cSyv3IO3Y5qL/a+iZaPEbUrzLJB4C+DNT8l8tPE8lKYnEhqb
PUhr8ivzK+8Lng3aSMsU7khA0cYtxDP1gZUlYU2bBTSBQnPtyg7WgSRYxmXhvoKBJS05KeQ4N3fm
qcMj581WVoAwsPSA8rcyWdFo5fYh5MYFQBCk6F5srDdJTHwIjf5DISzovrb3wfo632cSzluod0GK
E6V33WTZdODrLz39WEK0x002ze11MOGlj5VX2YTLAjJmoemo/YZSPe4iNDDzXbbXOZdan1agkWZD
RkUZPGBb9w+Pd12j0+S/mV86c1fxWIJ1VspPuGYngJYJcPsNtA+NBnXlgSkwXR6QVsT7Fbwz5l27
n9kwOrtIhD1qc7+G3n+KZ4CADE2qVS78EE4qioya2YLhuJAISyD1BLxlMYpYN4220jO9HKkfQI8A
2TTNYQ+KsIbagMduNL8WgN+B3GSkyp60OCXM6hxbYjbR7HmpUULspNLLkQeNNvHDvhqWfjzXrA03
l3GKF+v6c8/AICQd/BK261JXawLGasJd3ANefwY9+St/52n1aFCD2EqHuQyfO4+ESTFZ3xxTWajM
T1JsoAwLZ2il0fWwXvBBG/KPlByg9yX00YOcfY2sPEMzscnHmGnv1uPrAfynnaLvoAUDZkPI2qZ4
cE7SqxzDU/mWsuWQBjglDwaE6CM5qkVbKNa4jZXaCVJPsdAOJyXjLaO6eQFqNVN4ZwAvhODXCUPv
sfuQEiTYDlj1qrQpAni+BySplWr87WBeQb1APV6QOzEPPSHoUL8IaxgC8EyAilI8mTrCQ9CBiAN4
fXRgPX8V614h7EiNHZgJxYtxBXVxpMGfaoHE1W/M9ViWHbNvQuxFgUERsJ5JNWzltlQdIc/ZiPF7
cI5Jn9N53JF02RD4vpaIDlaoH4mbYtbiLwvmVi+/o2RN5+QXV9aDiGtvM7hO8D9ajSSTYdVLCTt1
xb/clQfVzUaUFfQoyF5DJ4yA6m+kEUz6Uyuwx/UwtCOvtM8z2KWrP/yYGequHBw9W86AYjeAg/I1
bLf7pkMus2hKUYa1C8PpHYF2rk+LSU8zaOrIJZHxU3D0qtIXy5gx4hPlsOoEDuKFm2PCu4wuUtGV
sz7kW50qrK0BVRjjHjdqBC/eJb+n/YmTp1suiiRxWFASj83VVrlNIkZmbVPWJfd3KEBRyl8Rfsbx
Hn/gs0LiTbDEFpI4ErYlh6Y584om5LnxkxvYVEnRUO0L5Y7pKJAkNEA7MJLDjDvvJuXpOTgtaWPH
1gMlJqsUtdc72rTHbuMOZEHAFb1q0Wx08zqV9x9UpD3MJNW9G6tIoNyrUrDFyocYDHXs9NdHJT1/
eEp8E05qOMonLeLg8RoPfdTiPLLnDQOsRT9F7hSqeUJm4ed/sbIO68g6VrYXCnVxDm402mvXv3jb
YSP/EJ4j6ezKy8sOJ0RwlNWr1/TYU4n1E3d9GPDbk2tpVnlvy8eH80d6+OFoJzjQilLAHDowd1Gl
WXrOSqyEajtGLsX2UDJbxYvmDu7JJLnz+Hw2WfUeLCVv0UI0cw36GrVRMjrAQRyv/0R9Kj1e/CzN
ueAvQ+GTsdU/GOM5+x3wQ1LM6AkVkxRP3lsyHqjjG5MtN0CsbF5XCfCeF/gLx3hfhJMc4RDcN0+M
tPrHgsY29RIWRFZyIQEb33vQkHBHlZPerR1AWqunAZM70/QCQ9i306DJU+rapAO4w1WK/qrtcfP1
zFSGOg/XPMzvXwAzbXD4+hFOpEonGUutmKj1OB+jBz0CKUCCoPxoA2NHzMBUgmusbWhvuVzFz3en
x7ofMrWWOnnGRya6MZfK9PgnhG9GN6JicLfxn9ksMA3vjCuj+adyHvJi3vzHC5d1zEIgGHCCXHg0
hurUtTzhpm1klr7xC9zW4D2dsbV1gOvY7Q2nQTZZ1eW5eX3LIZu8NmzZCEvG69mMVNYp7meJmaZ1
gxUhcQE0U2Kq+Zd3eJYmdTJ7oqkZwxGpOSFQSZe5SVBrSuypkwMBeJIDuHG/Z1Gxjvi3xO3jAOz8
gH8H/He9bFltwrmRhQ5JKPW752Oz0hVV4clKnQl2s89DaoR53XjGOH+aX/fFvN5N55ZOiSBmIYVN
BjneBNUMSJOCZj46mLNWjPK/C2U63R/Sav/lqNtozu0dfWWR/il28qdtfeaG2gXUevn31O+EGYMW
+qFgbPrOhJQad+/Wg1xrMe3Onuwr7Kt3GEa32MNMyfKmi2ghNTVrGRyoWg+nZxRyA42uWiGT2mD0
A/Cac73dC+MRoOhtpBPC09JAnNn7QHHHqDKEtJF2LwN5VuFCTbXVmVaNfckdWcOSFr1JynDUrirC
SP3MRtHq//nvcmrXxZg/6UaIHIDhmTs0w/vrQRrBBMMGKW7M6UR2x7I05z85HNUZfg1bOrkEMAlT
q5V6xN7ea4O/bxpCKbZH1ovDj/MJujD7ueRl195wsnlJzdi7HF824GIT5AaKX60+7wZBj5uQduIi
fR7Ti3t2NGkUxC3rQ1+SptEeEBuDdvJvz/zP3dEdxM4M58wrKhSMPWyl1YddNSwZguBg/kNAQxfX
qGJDPiYQnTO8Fl9LSu1Vqfhk8h/WgH7+d6Hq5JB62LoUodTHU0KN0md1PTSaZeEfUIou7bYjxIQW
HcYvkSYRMC1KrN9IEyL6wQWpCrW8a02I8ZKcxmts+fu+NLBsp26tWf+HUmPmhY78smQ4s0eaMaJ6
xUlwcPHtLExtFDcjNPQa4Mt50eFzwM0NoLvPzxPkm1HfnbFvx4E3nOdbY89haim06wCrMYmWgiCp
E3M0Rfwjl0bzthhFiUbzIlwATQd1GV8OI7E7ON5th3xjb4JZuZmEJKos2Ou0Zcq5XMlUjnmDjqeW
vQkk/geZGAFFjRWw9KHXk3JapG+iiXZcVdmTY0+cRkkCa/0qkUCgZs+ydd/hhnWdM0Y0s1yl+VWI
JieFO+YiNvphjOkmAabMlslw057VdbIDNhWwGUzQJAlJ8qiAgWkFUzLASWeGhR1BFqqI3x4gVDqJ
PLfIMlR330aCsfXRqrN5Ww/HvDoi7EPpjggK/Zo4INMkoV7NMyzGAIYhxQS4VutU23VQk8REhtsO
SQ386/p3oLxPP5BmHHMeOvmAE0wn3syyjZay1L/BPvQnRpr01SuqhiPdaUOZnohXrijRcdZ/79zD
c2rDzTZriG62UYnLI7TESVgmrmVFdgLMrpDTi4p2TpdO7UMFcL+gnTG4mlTS0kipj+IrOG4AL7L4
ichK9CFoUcAWlApGuqCs3vb1oUWVh3PSAjedqc4LJKgnuzYD8vMbLDI859qF8aYygXsZctwqnV/4
1sUwXUvEzRk+y7OVUqW+rUFer3+1RYo/RZ1TOiRXCHGtkZUKNpR43IqTG3oOeissnoLjwUifxXwd
kQGE55bDKlfs0XBtNLOlimBbkcDMDB5OIMpjo8HiFmU/irOZNt8F2/zHedQQjsIvyBGmoETggRXm
Evgwk/qbv1DKCS9+CZ4VDxMdXNS+fOWQhgSz2nffUPfFKOC5SxXhEbSz3KGmrngJtXYv02owJw4c
u/irme+T3DAEF/ocuT7xM2WW8zfXpl5FcAfEmAlZm9wmojg+liVdep7TCk9WU84tGlnzrPVzf/rO
Cpr44rRQ9HYcPfq3O/cbeNOphVDcwLMt+Tbacov5tR+q07tsTH6mjKRD0DAzw0Mj9TiQvvutvwxC
TTcJFKDGeco5ExupS1fQIcDdpMDRJ1ej4gTO/sGGhB4nFqG+5Te8mrL7LSrylnSk5lgZA/IXtgxV
jw4qnY5CsSfyE+HMYJc0PLSmUk523sg7qCz+zaTdo67jmHHC+aYqfp3Z9QQQhkyTwXkIn2N2dSpQ
2qTEKogiz/mqr74jFtxsYJ7ngBaUPfkDJFeIYYGz0Fe1TofhU8hKL4gkcu0txFMQZUj6o8scVEWb
05WEXCz7fmbl7PXANL2QwC6kmPvRO+jjD678aj50UFrl/aksIw+KDnvwTu/98MNqXSVkDUCFQ0Ef
sm911Y3ybVMAoKNMAZeWcZP/23wlJBG78GCVytpSq4QTjHDVSWCyBYtJz9ngi9g40ZMtmZ8Nbi4E
L04SXar4W/hk3/3AOxjIf8eXM++rCyAtjwYStfSK3oKV9QhGkQYCsYB0XJDazFPwllRLKB0rSeEh
4YtrYR287jysZMYSPGl9pvFoOWnvP0FrzOHqr+zPIiySw+eT1KmjZSma8PXlxeGg2EID7jmC1wBC
WFM/sVkCl92OXQMOcerJH9gYW/VMykjelen4bkdIM39wOIBnsRg7rfKVpCZ6teZb5477b855qup/
1GAYU5vvDzTyvjATQvc8RjRXb8q7ateJbaJhKnCps8DeaRnuVuQl7Pz9aGgG/l4Oj+UPCJfVoa/t
qfr0iNSGU147YLMkDzn89rfBqUp4+xL+dVcpRRC7fVic4/n3t/2veOFtQmh00n0MyaeALLXm2Jt0
fbTBSnszvpygbk79ZGOp1jfHUt7nzmdidlzCvKnA9oSW7eiTZA33zW4G8v2uG+dcGwZlyH6SMO6c
Ry27MNiYFo3nPBQxd2seSTnc09UoFI28IEz5SuE8VUox23x/Dnq9Aw1mk6ifiKbbDyZGNoPqB5aS
CCQEsnwdgs4rT9Vv0QmJxqc0rWFo1U16DKsR/LemT/mZmTS5FUfqoT8GsXPVRdm8En/lkVZ3dJy6
iO+h7xJZ+7ajtoOFszzwCzV3Veao9rG/pn9gF0mugx6l/UAPtvQ5qE9P5shdurRMh9RB2SY722d/
HN8NF2x9auWTPVPaxlNVtJdN04Wp4wV5ap3Xd03DWRqOffYpDhc4Co+QPO6LKHCP7dKj2rHgBGgC
VHvhFfdS8Zrb73Rx+21k2Q2cEBb0JHFPKyhrg/4yZwDJ4NE9LSeWFhGKl+quICC7E2o35t/iew2k
yja/zRSaRPjInxCA5bHXn32fHlxrZflUKmBUgGOVm3kZvfsEQtOjGQhGc+apu2ZfisNGN8nXvoF4
UDnjHtvo1nQd0XcC5si67K0elOn7KHxQDvWZxhonR8nNRPPhsfbH3ok+6QmqapVZAnF40v0toKS5
gDKT9oKbe9WLRSijB1z7QMGzS8QimEHBy4tK2F0KI+bbZ5+J13PKD3EZyvOssCWxQWEY0eB5fMcn
sjJcAQM2ZhTdFzb6nZh3TyBC0xISWSUvzHnAAmdEVyzplXtY0LVqWHgBDrLKdYlk6/p9zMJy/x0X
gC3JbqdNF+eod7mul1c61jf8vz5Jtsk04PGELoo/FEc+7uX4osskbSVLVpQhW/0N7GPHw11wXLkV
Hiz6abAX6Yqe3IskLPJUf28Cahm8THy3TzlTfoQbDMnBvVcWbJh9km2lBD009w90IfGs9sOEUXCX
B7n0zXZfa+dJou5z3sfAgTi3cKj0GWJaVY7loBDQ+VkibTPBXhnqAlC7sIUlDl7AHg6GCWlchQ6e
5PzTqxAbX14ayWHswyH79gZh7sJgH2ZIiwnW4+TaWa9jUGVP8FhKQjovB14Su7doaH1Xpa7NxsCy
HW3XjvNs0H5awXznc4pBnpJMCKzcAmg7WnVGCvMzmM0kJscFnif6K9TFUZ87PDP21+KPc+gV66cY
5CP6Q5sTl91u3e9CjWsl6oanJ4A050R+cQLI/lCVIr/MZjEOij3z4W6JuAqqXDLATZUoMTB7way5
c4HUdIMHYVwCLrNmfMd3rfAh3xTEkuYpjQFDFeyrXKljdu0UfvJko0iicYRj+Yq7jKfAcYcoBOns
0fmg0rluvHnJ6TTg0N4Jgpa/H3yUTckxKmY58gxcx0qXwM1rlJB7rgHgLP/2m8FI15LBTEjRqkP1
t+tnF40xap9zCdKyiKJbHGEHIdxiQtaoQHYdnbgm/l2bva/ZHsrRMEh8QAa4TxMnD/2TkMflVs2Z
y9oKQhhjWzcsGFt/mV8oELt0k9P3E8pq8roiK6xhNKnTwzTIna0VwV6WUDDiykbh4Td+/WTXl4pu
bwJ6GpB6IkyKl3bVN6b5efjkr2ifw4U5d7qATMh3hh3i2aj946O4NIVyrc+m9aJ+9o2AJIzAYD20
Gqj/uocff77KL5EQ/s+ilo9NWfmrAUslC2wjA0lLyFcqb2SmSENolIeERhhL2yevXJjX6tqLciWc
jdaJIhQFBBwfsa8YVtOzVKwWBT8aEQWX3Sy5RZuVSQqt/kt3Gio62R8caQiu99LL6rK5l4F151s2
P77ZSdyJGYBcKkvTJtbOMt+5lOxZ4HasJjpPqpH2IiuRnyvGzD4LFxv3b0X/96WW7DFC0eMTQNG7
NH7z1PYU+kz3DcBIK2guJ9Evq0nkNsX6WNz8945xjKYWbBtUOexEQrCzS4KcSER0J0Q1KDiq9ALW
TEekVLROcFZJkDXXwizTOFEYiUOqnGFTHoXWPZVtC7omwX9cPuv6aRPP1KhAPn72az6Zi5845Sn6
5WrtFQLlRhOIH+VBF56Mxk10Xald/fEduwyks4tgXyMj8V1pVCQy/VX4vjxCHY/UyShM82c1dcmC
FB4bmUNH0ewYgFdRUNGwxMM1K9q+Q3uqODgr3fsoX89qKtTO5AT/XFhp91xJwoz41e28hMMs1q+y
hAMNYcVDK3FGrK5x+FHYt+QuRXriJDis3NElrQ39F6JHQtvnu28QZIfnLQTKZROnBikBGqtP3egG
9mZ3WYJWY1oCTyO3PpBeVwp8TpwPXWJdD74Nn6p08s1Kp3yOHK5330EbXV323CyCV3phaoDc/P7m
MFD+fNWNEscmcNrVlIWhGwwARLaGvaqnnqCOqcfoBkF02vtISFrc03jyr8YP4pzhi9LOoVQk9YL/
PxBxn+g5Gi+bXcDWOkwvNoJvymNpeiWrSVgJ7Pzgi5xJ4hPZOseAiCMmtDCV4BGFX+2snO17OORy
i4SBlFK0G4+mxxWyDVpSegnqpK/VHAwrgiMPUC4pQjYoPfWZBlYxFz6GhkK+1yBPJZjznNiex3U2
+OF7tx3VI8Die1ySDxivYTtkPtcuVbU5CC0CtgbUxAgChvJhoQDalthqAGcrBSLNMOtL8Oy4HabD
FGevdkwZqrXHXCJH9zasPxqJpooaLL+51nU72CM2AChiDxu+BXGjhHRuSn2SE16EtKgLla9NEhFs
2jse9Li/9o5s8zm7HpUFmNRWOAoNwN10a75XC7Wi0HxWlqdkKknOv8B618s67BnolIhG4c2QakfM
V9szGO1OPeK6Awj3twpgdcI4h/GkiF+jsrEzq3CNyqFv7KG9gWRJ9popeM7jwVrJ0+RYVRoPQYel
nc/x7prTY/xsBDkR+sAXCm5A5YUsxkug3td/Vrv8P/DeWsnT5qrj+2yaZBswxQCktkd9R8WkFZfk
blkfRSw7yUCS8zSfVHVKbFfi6K43SikfiFbGiQHkTRdvgOQZwRTg9OhD3KT4HxzaLX3ZMcPPXFhX
5Wa1Do3ITq8bEw0HhRbT8OJvb85g/QtU01tIQGsplIH2GS5B4kaE6e+zPushcdDwj0UjD/u9JeCf
fNmoMteTCXpYb3gavALvUxzfYHS8itMUxH4j2nW3S8DkZJLN/1oWPhDVRdHutjQhnui7tQPcs99H
B/urWYOJLeLJ63E9LT8PuZcGKExyD46P4dFvInUnFhPu1CwfPqJnRGMHsjSnA85KrLQxj+bQCnfk
hx1AK3qoSn1Fd93F2LyLoMyCgdNvGcIOrxymA3+bpcfY3SWlmmiYk7/YADb5dKZuiKWVS4cn4x8F
wQgLSRGi2hm1nEXS4Ti4Ppnd742Wa7OwjCIaT8MiCaBR/abz2OCh0ooBkk4tSNEaFr5H70EZZsTq
Ue3oGHIs5E2Ueul6A6LfEZppAu4pCuMCkcLUOKM4rFLgdzTg6fNByhYGnGM37AfiUGaYs6NP5H5B
GIwTuT1zZJtp9+TA1uAVULiZ2057FnepCjaQkiYFnl+VqiPKAjvyrqZJgKAGvIbajMyMkRfd0FOZ
mhE/2s01XaZBuEgO3l7GqO3DutGti5QwL4MumiSzkCZfAacUBOhodvNn6v8RpvnBQk1Vsn1GI8t3
qK/Q33QMREiiaoV+kR/XYSfJed3AnojagcIf4QazgZL6cIb5tVyysP0+Hq4u3i9uqIBe0NV6EJw9
J01CaKpc5QH3lbeeHpllADxrIkxLW/+3ez/qHMWRalEdfOdCc0TGe4tF510sESVN52Vr/UeDLB3G
1ESyTEJsAy7CNlwjo/parmjekxvvT4dCAuACq7mmKXng8zMmy/ens5covUysWQ+j7J+5TqDck8+i
FMzff4F72404TiB3rRTCDjGQf55hlNL8zomIWsUBWK8dCLHl63IrSz7f4gCaIAy0A5cPYlDQDUGq
lz2cJO/tV8Ewo4EihZI+mHNE4Lf2Xj7W6i5mz24IP1+NIDw+mlBtIlZfeNsXc0g9mtwm2Ts6A0s5
DjQNDNwdpyC4BbeYvmdj9TqCDZFRF1WK3z4+ZjWyYvW7Kdxl93cVmFm0Hj/SBL5wrZ6ObQKjz6ho
si3jTNlwxxDk5/s224qXGV9ZWZCd/uYFcBodR4nol8/44w3udGf/J2wXmpcdk6FYJFrj392nqaGL
TS0isyjrYgWArQ5IThEfT8x9YY0BCvx4IqoSEaz4gxnp0fl9iLQuXsj9V5uczInTrWdV+4M0wlgV
uTRTzmEqJcXUX9kMI+YH6FwywbazcwHyO6wusPog/nBpD9g4xA//2cFw6hzYuEfLFMZHWu6O3Ena
xK1oKieEfZj0xmwLn5hv1ozJTNKwIuySY1jU4wJYaBOXoYgnIFZPnhdMYLj4xvFi5fNWURMphJYX
AVfA+gmEbHq0KuqHSW1cSThTEFFC2fQ+d+EbO59JIO0HzXzULJqmzZDkJ4sJIdMMw4yz1TVO04qR
zV4HUWB3Vy0ib/uj03yKYnifGYrRlntTGzONFi2WnFfmg/2ZgbfOI9FoK0qDGwBlc2Kccbtq1IuJ
c7R30iiZvhRjB3vXzt9KCK32ZlrHj97kJ4M+BikYXAjaChq/a1cu8NEugfxZXDxt010OAcsWI8jG
L/Qeg2XKTdtABjii1pPVUr/u1pQbBEChM4yXuVEVrFOnksetDREaJW0VSGG5G2zG1SlEWSaFu6TP
D2dTzw7zAOyxu0YmNKAUa23BcVjH5BwVjjdCtQEQDPNF9CAl6nyYLlBdJM+3TJ+xQGh3ZtYcQCAD
Z9e6gL7RYSm/TZ8SOEceTLe227ywFBavFxXxHfEXMgXOEUahMaYk+KxHO82vcdmM4HLfU7eg969v
c0KiEQZL94FSzdX7//BKLLuSPhmKJlhbsnsYFVt0ga6X2w++abl3Gso8Uj9IMpISItvLak3OieH9
t4ZP0IUvsNdLBoV1Eidlp+qCGoWF11wblZyXSVnHENkeMRMm6QckitGEjDNqWSSRxnIcWmoQRIa8
d78hN87iqmseNIMnm58WyY+QHguFLcQ1WUklDPjabN6pWoJ0pezwBJ4OGCocJrs+JuYngTOsKWnM
/dq0o7QJJVmm0gj8lTXnYwU9rO9ATYrTmCaHcsVz1IAgqGbqS79jhYdtlc/tWvn5E57iOKEfA0yv
CX/4+xasMb40IzoE4B9gow36ZIiku5E5w1NCEBOokfn1oW7hUEEIxOthEJo9vbhxptLzM6JR0vgM
Z+uBpDVKUc1TWMfmLEGUC6v0MAhimaAEKWUt08xF4nnozBc1ReiBrjIDrrrEJoJ2PYY9Ems2s+lR
2/+QoN6qWmGPKchArhNHHev7po085G3E0u6fMFS/EH6lxqLNIVTLBKiH0/U+qJnE6nQSWxNOJp3W
ad7uSRi0i5eqacyWhiBzgjrZ5DLS7Fx4oZNpfCtMRCvMCzbwrkjaSbcVKGxSPJac5378tBrVwX4Z
pu1V738mSBqX2bubIlHiksGJ4NvcqtJW7xLaqcclp7S6fWX2ZOSWHnHZ2ALmdQF+42zQ3vIcgkZK
MfCk6PrrxQfl2gzXGVCQoGlPnUiQG5NlU9a+u52FaJV7DzHZbqGI7rY7/osprQ3CGVcOMOe5A/uY
yZs0FE2ARmu5Jp3iNUUugCtzaq0uWcSvUPWh/77qj8rQIBNVU3/Ttsh16tYRtGIoYRFAWZvAEEGw
kxaFyf8hA/yYO/CcGTuOhg88fE6KvDht4uzxTsXGGcZKu8hBSSjFHft4Phi57f/SNsg677ODc9JC
EyMpRsyeKWfh8XZEdj+dJ6ULKLMYnWDPZ45S2XzbbF265MzOGs7NyV2Z+9iLbeDzwWxwi2Av90xP
PAlou6Wvg4DRgCrNZY0as+i/gHQu9Wn3MN3xRUKrtbGTSaRhx5UbafAoiIiab3jri1LTR27LBCqG
Fl8HfHwZLiY65dnBjpYTTteUdCFG/FEaO8Y4xGkQnSquTWUkjub0qbXmj99AGzp8J9zVlQbFywTQ
d+VKvhfhLi8RhmAhmeEiyhxrY2V9vOfFks6+7yOm9f7wk/S2M6ipcpXYPz6uFRy9nQZurtfYLsVg
WogNo69ZSsF9Mjry8ZQ0j+5znB6TdJndFfmOb+9HcM6E7jBrnTFQe9nbH8CgXSRprdjIYGRIjdTW
0gKQK6g4Ac8jVahPUGCp3IUh2lVdFiVMobG9d/InMXgYd0WL3MoxmJNTyQmmTuQt9pRxtnC67WG8
08ywvc8LJ4EjH3pMlrhgwKoZxdS7qQvJSaWam2qV52eKqRiVcSaGEOCxh1auw5OIXyAaMgdKy9Gq
NhTRxf3DLVlA1QjwplGzYi2vVXoR3O0InZ74drxPVVFIJzd7Q/pMEqLaCM/olv3gMary5DpFpUAg
26wJEImhRNvMv+5f5B3RM41JLem7O2AAAI4sDtJslrD7QMoCVJzQtAxY0dRyYypxPW+I0FRIgFlw
KQ3OtT+dDv5IctIhWMXjJpkU+9SGzew1J5kCdOvBvh8eQ+tzh91qFqY9TpplkRgXIVsacRJH+iPR
OfGkJL704aWdBljKoLabwnAMENrEubPvVYVonZdH47eUdem6KYJwa8SIukBL6ny2HlUIweMHQQn0
25peId8amaPPn5UxkbWD8ZIfH6thAYdl8glLR50Of+d6hosOXYAodKlW4XVGWRy7h1EI6eg1vZki
ID8xoM39RFxCkXnlMQXAD3vGVOAArTnl2huMHWutoAA4WuewcgJemX1sDGFRMXFk5/M/Euxw3iy7
bNAVyvL3bv3BiBKf+t3gLhBEp5FGoJmrRRr9y9hykhK+uhfK/6QpbjzPUglUwg6uzENhl3K5RIPW
WzjJcgdtInfjhpZ5R1YUfvzBH1BgLwoNVfuPMAkk4wyrqvaO2ho8oUOy3hd78eKZYty78eD8Jr6Z
sBj1+Ll6IoaLENNd9zkm818je4/ftwZ8P9MnI6JLFqTSOenJTyUnYGpvoZX2JpOBaxrCbZXX+k+m
Ay5egBTw4fI15M8nYBZ8vXJ5/v9G0g293E37qbOgCvG5/V1dYVQWUMva11gCU4/WLVmgEiD67S88
z0gHJSJfG6n9plJMMrhlFQqP/CmicsyiU3sR9PYsclsbtZqAieZLvpaY5cm5Ujib8yeZYIGAu8xM
U4a4Net9xjVxVwaUkS7jTOF2k0XSthAy8H0Ng57Y8vOW5pYn0UCq/I/MAsDWT2nQzvtxCJrrGC7X
C6/ZAZs+v8vMNvlStw+IK1o8NWgQn67JubLKnmbGS3z5HCBJJRV1RKYjZFUAoLDNG6GZVPnhsUkr
UMl8gTbQaoVDEd87UApnmtIZVQyPlrr1CW8gwmKSnW4lk2Fdh2wJUVzvMn1cF3Hp9UgM/Lnm/4YQ
tIXgzY2WkO2RLEXen3qJ5AtlA+uKlB9CRwZdOX13m2AGTONSvTf2HSnlNF28Qw1LE69aIeGWYZBD
xHstvwVWHhPQLavxvlWL0hDI8RyjK1sg8/VcIRGp3K5Sjaro52bKpL36bnq36fXiW5tfxwYEZ8ku
J1wCpUiZiNVcmwpOA7msNz+gwKN9d55rV7FATn23xdnKPJsDXIFmjYGa3A/KkSJ2p+Ar9BWGibot
IpwbsPTA785QhXBxJ0bWc+z0o/FDUrDnMd75s9ebs3vw0Tf7AM2hDM5bcJoREVQ5fmS0eTg3zW1X
Ke13KV8sBEYMyU+g2BbMPmeekl9QV+PBUlW5yfKR7YHvpNyKKt0N6ojxY0v67TcqLArO1gie5xPR
z1OakwcLOUOaJhu/aADBvaKMfqC3yLIWvn++BRt2z2yQEbSHpUxAJ7vI8MSQimcSz9n9M5CmRrE1
nJH2WeHrDvZLLroJ64F/6sV9O+nIU8Cx/oK1sZdECSXLWikTXvHZKPfpscN7tKztevhGJKxsvpuU
IcT5NNtmh00YSp2aSMr8OW5+LloPsMN2joN9niYXFtH56Tx2NicYnpdpO1Y/e2+gR3pWIlhU5Kx6
EhAGt65//hDBgCAn6zzL8wzslPRoU4u0LI+ONghXL/uMzkCmcF1BDqnaNvKx4z/D5CLerLLYanNz
8iw0XMaon9UrfZK3U0Bx+d5X1eNqaHSv/B+ajCYVjx8K37Uff2aMEB1YmJXtT08iUr8aOVyFpLzb
lwXtOgUgha/MBxmdjA5tkS0YT8T98hTV9SVmL/9q5aofxBxL7T1+liyIrXRz4OFhdBTGvYJ3UaX0
jItSZjXth5eIbGX/7sm7hKFZaVmdvZuhg/DesUmUZkpCRhnmDxjtKnTkGN+jCiHmdnw6lZ3B9+jW
s1jgcJHlNFdGAW38zhc0pKdFyAERMJYlzJmxP7aYl7K6KuxdDXMaD1FfDeLyfP08Qw7oa9yodLBo
6nXkWgz0+o3J6Icwsurks3P/Hz+uAMZMjnSV/HD6KQG8ngcVeqLx3NbcSXRaSRNZVm5hE0xgcqBw
ZaRp91YsCZWtWpfSOnNAVQ+4Z+NkvaNShWj7WPYC+1XnxukZ2WEb65PMyBdByV1qisPen1wCZLsj
PfATG0T45+nAsve006sd0kROacfKh93LPQsqI915fRYe3beQOCeL37FNc0Kx2lpHU3EL6GX6Hqrh
/CJjehs0MK4dpiGA+1Wm9KbfYhjgoMMer8C/qX05qcCkQjD1FRNZYFGFns0nt7+jfiW2AlZ9obLU
CYwVTpg9Urx86E/NgIVJG5dstLqhI72bjifAI/O6Qrjk1zGvvcGmYy42gLBHqVL8ISWH5TlgvN58
kSHStgxUzIRJL5SXOmNqUtD3rsY+0gieRHerBFD+ZhJ8HBZh+B4o0Kdqfxk9v93BCBjmOgXyDVaZ
E7GE3nnkaSbyvr8EWsS/m7hYHtmp3pdEtGle179jsW0UxcxA5rwtfEagLQTNcQTfcpp43+sh+TBb
DICA+BBFI25VAgs1zSivSjTH/79VXtr0ihPUSKHrK1CC6pDK0bM2MHh6PBq4yN4qO8eOWarw035c
b5Wzm/8qlyKMFWnSYxSx8lm0gQ5Lp8gm3qElWSqhPAk7e7eiSRSx9GHpfKtT15qMPgIxHo6+zaY6
eVdI4i+1JUs9Mc/xiWuMjikqWJGfxgV0p7JlF+IxAKbaaT5xdpwifCnrqxu5DxxklRWQAPOWHW+S
uVe0IAA1YheIdEplwK/ZyK4K/W7Cpj1jn809ykVDi3OkEgAXPsEWzI+vZoun4nFuVjyf6ugWZkHy
HXXDHmICjXBX45qQC6zCS1s4b0j7KTm/TJ4j4h1Gfz/RwBZe4GP+U5SK1XjIJVRQRQumlHf+xACc
EqlYpkMiFwVbVe18whiWW4yqXQObUCEYqyRpUPLCXMrdNt6uUNUftrAPq8w83bBNzmVUxU3M2o3j
YttpH2tD/YewHgHH7M+KWTvhfxn6b/PX1ddqbr9keGSsHIQEZAu+Im4k0x/sOicKWFNExi1gnE2R
Ni890gd9orpZ9musQ011mDPcgEYu0aSjbRP8arKQLsfpm2xkL81dkjZ9oG9vviyazhkno/I7tJsV
cIeHVpfGxRbac8i1AHNbrPu8/sc74rBt5Fjgbp7lSDi5BgxGOVU+M8JrmX/pQhywYS8QP0mfOu0X
KCYL9l/xmneeN0YFsuXMVafTHbU6ePZuCSE3/GVyC/IPKS5r+DWmgmbwEfV6i50eUw3ILgTkmm6U
O4vKys+zs6/RsSmlVwK9Cb84j0cSwW8eUUOc+dvNlatTt7LUs37P/R1azqrH4LQvkH4FcpqRlbrh
cGhZrNsArgpuQ4L8k9p/xuCX9ErnWvPjSSA8y3u7laBEu3VHL6OaTz/YGrZZUFPJKhGzS3WLpo8f
TwR3wyBVZEuUcUdYoXiVrra4/dQPjFmRRROBSR5/TF0cEo+oVvp64XAWbueAt7yJlbXUis0BpOia
bJ/a1KHmmEUcgFARSoevl8uMdH+g6dMNVFwk9TvCf0C+/dVATWwJBgP63tvkFEtFJCys1kX6js6e
9mPEyOdAlxBgRi8D5031hfAgAWaXTKEiudOC7uagmO3wzXIIXxvwyDobn6yfp8SZz/+4zY45P0k1
SwreigtVfXwXuy08HM8iVZMAPjYTseX6fy0KmxzSi7ghvEq7OjwxrG9QFDuxKX4u04t0a2piHc2d
LMnXyH/JlKdIqnK5eNMCvOmvLk0HJ3ocEKH2rYjrBEzpMJ7h0G/7A6WOusQAgs87mQ9JbG+72HyL
kqQLjiE4oUX/isyPWhs7ExVwnak8qHDc9cTCxO+p5p01TWiL9+pWf3ZPU6y3FDNuOKNMjwRu+1Ht
JWZZ6KYJCk2oV26vLwhOeHUemehHwyrmAoa5cLagOLX4LpyTrZg42m494cFfQqbDb3rQ++mcbaDQ
J7rrPhfuR5dTKp7wB5XdVcFO/o1TFEzQJxpyCW2gSFVAaWGRqD9+61yuo1ppOzknvkA8EUZaWkZ0
/lolyqlzAquOWYgC0fLnQkuQXHa0TT/EQ8Y9E7719tJ33wzNkImYlJTF1rrmIykhTVJR0cYz2uq/
iB4h6Ye/Ug5X0Q0YTMbQ1u3yA48xowfKLBzJUhml6J4JDuO5iZ5Uh4q5NikQwQTxBC8RsECqiW87
8Q3Y5paNhEr0nX7u3FoKN8kpcdUSsMMw/KVEGi5Y6sE6vddKnnHPj1Y3HiAYk/Di2O4qJH95dLHK
/iIHDlDJHWF2FKCJEJvCz8Xa6KwJzs/F5Il9kedvG45ayA6A44ncNYMPN6gEMxaTi183PyQWVEjv
RxkVVqOXLcsYq75wK147t8hsUe/uRqS+XTPmbAVuKc5s4d7NMu16Yg3tSYF1fEWA7hAmz5MNU0Vc
F4OhokifnolyTNgyGry3MATZJ8WTlSTS+Zyq0ay0xZ4UsZh++5D5qxx4MDbLw92IhNI4yNAxJyIG
AgsTIl4JcLCvHqFyWKGcRMr+18nWZkQ5Y7dtdxQWPBYwGY4wZ5OYTKYFQyZI8n+SfoxRK83roXNW
fy9wO95FKYyhNd+2QS7sCPJnHcCyEE9POIspbucz/s+kxyCvpi9AL9fF7tUSSzDk5t/w44O5IXEH
mtpoRIikHf9lx9jXB9InNktrkcXamJ95CzMWhFiCuqvttyfHtWPGxBLESHsYQFc43gVM3E3Lq9U2
SHn85Lqb70QJjfkOayUb7nrHDsYypKosBiZxJedbpjsg6LVB67escpQ9YGl9OcyRQ/UfD/SBqu3U
mHwG67R/IEiOhpKxODVl45dphQold513JiMiACOJbtmJ3Q2dHlmxhiPU5Jvq7gRzWLkklgcm2mGU
JzvcBIZGZ8ArZ4XzoJTIjWVU3YSRqaavtBaTzYZLfMELy7jdV/YfAhSIwDdybk1nW+BrrUI+/k6n
WvPhvjdbxWB4vt1+6yTKaYbZZZMAywkB4Km+GmOAdYNNSsNZkm8cjLEmC0KJ3Bj6YxQYJNBFgBlr
Ff3/ha+7ZimiRww1NirqQ8juKkZYJ0In28hWlelwehMSusFquVjDxnqs4I1K10Qx/u9THtFwF3s3
XNWgRcGtPqN+1NKmhLq8Go8NuwO7GEKKg5Gm2IUFsN3oCSVG7nzBcMS3j62jPmKwiaZCwAINDCE6
Nejl72x+8FU9SojRyNjd2PM/4w2Sn+PTeprvNgCHVJCjYroicgL9gc/cnPnT2go6x+PL5DjS2Rex
J1m/wEY5e3mrVRA9qGVP3SVm/P4MrLtJA130SvMQCSVKmUKTFe8uWlyVuGeh7H1bRIZjhv0p33Vo
hZsttwCQgfzAyugv+BLDZkmrc5ltJhs7ETylSw1x1xGmDyYCOu+WdzU3kNT67qe9NpV2/KxhX9/T
1OcWvj6ItpMagt3xA5pf+74UsCem9B5jvPkqgThWxPT84iyxvC8VAj2jX8iYCdnFLQpL7QRy9Tmm
MNR6Rcq4NO6DasdKwP3NHxY65UD6mrBHsTW5gZ9Buk6iPb7Z7+9JWI8262eIK40glYm9/zmJPPJA
+iVXW13JASGB5oJQc4caRuhBYO3nYR2iVJwdXvx+YovE75Uj64EnYehM0N/x6RqITgk8mlTX8EvN
CnaW0Cy/T99MM7EXmOCEvwc1X8u2sg4ki3XAHk4MWhiOW4qsecJ6Cbl7XGG2mHVjFI/FJbhSLRRc
VYuPDqsGTB3fH4RGszUgokJRtBQinE4WBvygOgCnzbffcMNPeVghm0fy70fCvHgMBOkSW/EgaXfP
6NGSJZXvTn8Mho7ElM8RhYymQVVZvjh5da8om0gPZwJJ1w0KqFnuKTLQkgEMLX3Vk6cU+KN+C7Af
cYbMuprDuCPE8EeUWuOs7jUJUE4WF/r29JiWh/DGwFOGLc2EokMxNGvbscxQwOHw8HSRbGdO7jjp
3GaHt+JeGSicB5a6/QeJIhJuniKbjzODHMFUjNLeLWFYi4rOBBdxYDbQ7SxhhRmlUtAqPllRfwQl
IeOgDDE/btyuGn7aqE8lXLwEfsUGbcy/N0pnbSZ0SM4j/wvgRlWozDSswhx1RRplJb/UJsR/98fa
ZY9RLU6H2jZE+tOrE5ppjHe4bfhuF1iRPrp9ROuvqiRiTBvPDOAqXW1XYQ08fRsD5nPcH79UKIoe
HR3fKb3Z6bZ7nM+YyVzbXstLpkYRroxkr+Jc0ndLF1R7Fx26TWAAGbt3Ew5oYqZqKNLN+pVTN7gh
d6Ykuc9X0DPG6543Ny326/cf07j9ePzS4rhZ5K+2F16Plwy4C1RPWVicJefRS9KS1EFjapTHG1Pu
qJr2VXVj46ktS5PNb+Y83Uc8ZeZD2kuIzrFKALeHk58MoYCVqpRFzj9u6hwF3OLDMgRmBa8qkTBk
JFCMbbTGCdLKlnMERtsNZl05W4iAgHZPkD4DDCtEbdWuI8DTComoI+CHmhZqOCM721RADrVZiSAj
/tVAjfuXkdYj1N1xKwBJmBbK4uL2eXOoi3ALVoRF88oFrZHs694ISrFRtRqlXwq2pm5NYWybQtf+
FivQR93NOMWnwPCTJ95X+lmlMsY+qLnY+1FgjhWGvBopYabZ71TzG0UNWZSOi1/qNKsA6zlPqJ19
2U9vu3BdVPSk4oCWGeFW3M3dKTRqg1EgJMYLcjWUhyIvb9FfW8XcYwmwSB0ibGS6Zc6C+5Gt3w+Z
K2C9h6nPyY9qAUAJs9P+IdGXgGMipJB24X033FwRoM7+ThtiGk9u/TYpMBxNyDrFKpVBinzVawyM
sYDt0DTjhKbDNJ3sGDhwCxb1+ZomLjuwso4nuqveZIAODDsezHlncLyPxZ41gmFiAPVgF70q07h+
WLCkwl5aP9bmWyGqcBJR+mpOuvTUC26vD3v0jm3Odp8YxHbOclPox0wujKHV0mAsH1zkkRxyWgyA
U4kvDh3CCLtz3FmTCKNRqiVfJmfeiQXT9+Zx1yRSBL+t9W7lEgAI5STJWjx9uw1JDYvrQj6rcmwq
ag1eFU3nEKsEa98xR8A63j3xi8Tlh+KaBpkWITnTCYYQUDjCf0FBmkaGhrxEddCg4ss17oJXvQ7l
1poER+VloOz65bNuYeGpfRR5ytgWAgNquvMcqIvkVsX/enX+vlvqhMsuAQdO9vjDqn2amovqPw78
0pN16obEXFGyeobC7cyMNixhm/czaL4MiJ12PeQYYKA196JpHoj6zi6T5iZMWSMKv81fpZ9aCFrk
hXE1AQukViRcasrl5JgJyBjHD1iiKuVrS60DM1AhK+GHDIbE1JnBdFMD2RK2vjyZFFnFSWV0Z4pm
KjP2WufPpKs5caweizI5qp6x1fADaI8aEgGZ4DG1Wlaszx7by2SE7U908NERo7ZzjdA5B/knmj3K
MFdp6qVm2wMT85rfMZvDMAgVDqCNex9jmGdGBOfDZpXdFO6hfw/bD5E8V9mODiAoXkHMh8ZJyTMv
y5XZcqLLmYdftdsy3JZgG08M1SibykBM5KO495HW4zdpcVbNKbJtaU9Zebqevd6jb/lQ5905Pf60
ZmWQEn/LlsxmrHc3xu6nWdqt42tnW+wbXzWL+h6kSP6DKkLeKE3XABMbAMcLcSE6VUZvx/OjNqfi
Xkmu+p4WRjrNPd9U06YIq5bKF9CN6cf/f2SNnxWJY7Jxo2I/bhVUJ0tposBnHuw9CEaZBdM5/7DV
MlL0DdVtwo7HxpsMbPS01Cb9RIABm56oJN60SJ8ggBFAAKP2v65vmUAYAYpYIyLBtIWXJ+U7bWlJ
+rv82e9eIVVSoGSw4MSK9a9TdRsVaXsmb62UcIVtFs7niUeuxb+RWUhpvoT5xSKDYAdzjznaG9hD
hIhuSUCEpSaeu/iT66Yq0DRbyndkHsWkVeJTq3dQBsvhwYVml5MWsxMtZhMWg4seTiGq02kLtm3S
xw69QxZkkw5xljrQ8UdRq6tUR0eNwuAUleKkpTqO/eZxiue2UWW3FfdLVKGS7WJPYeWk/GOamUvP
G+kUrvOqWQvEGXkqr5Vs260d4r2sLkzPmYgFl0De2h53m3fhKK7txub2qUb7sZWr7OGvGCfJOPn6
NzPJjy22JhvImqwNVBEFZEIUsBLzeo5xRaEWCC4UM3KegWq0MEqUoerITfQC8dh3PnGepHSmTUoR
X3+c2TR6NkD7wqh3yihnDGGyl49VVaYn9cGvt5rg/0fqHt3w4AbgF/3mMJyvtMQAa0Pbk3xCaeVM
+godLiURuTZwFX+IOH4bnhnh5xGt5v9ysKcTlF5CKydmCjZJedvga3KQ0MSDHs69PlIEu1D3OYld
bh1V8BqKMv8uIdt4WC477pd//fHix+TWShao8wPvAbQ9p/XOI8VcRk7S5B1qAHh77EZH5/+PLJRB
PBZuo6lv5Zil12AyfHZoTLxEFfTQXklWlfE1VZYg1QhPGF9WdYZ8Nnw+mreNXGSPprP1o2ZyyvBF
LMWD8rJnlgvn/mhkOEwqUtBSo3KHQRH55DKvw3u0rl/3O69Gx8xTen8ZPXPPpB5yTGOUD+7ehW1T
rJ9FhkVo6weyHZvtfYMIwlzNEanOC/+QpFkSlKaNyeRPQmIwMh9iv8fjtQc2/kzy75mzn/g2TYQL
LKEsYkCMkdygRLMF/9AnOo7gcJwmkrxfATDOGadSDo0JZFt6ItAMgTMU/+5z10wZzAVR433Gycm7
gYv6e1Q9vNFmLiggC9g4OCRMmascdOs1Is+wq7CuFxDSCfi8n6qXu+hLg5hL2sJmr6pHRzEBBlx3
CjZ3GGkel8xAekoT5RKrCKfWHfxVokfah32pjO0/WdpxmQK7x9iWkZSlZ4oGfHFDaZWlYr/ufeJy
SXrF/O8K+74NdkudNI7QEKxa/zoKKrK6lAla9Q1keOawrRETX2dH8rThQRE5k570+r8feLh0JXn5
VsJFDJ91kA0ie5jXO67ipvNLkkg3QZ4AjK9XHOrejW/e6l8Io6DZfvHWvCIY2gMGr4YrDNrCO0xu
s2WBAUxBtDP/bbKpaX0/cDVh2iYEDBfhWPva31sy0ctFzV3FAVaoLGW8O7Ti9KR8C5UnrSRxZEzi
J/Sh2VVQ4WzF3YYXrVShoc83mQSWvyQo0VFcdGW5mNY4Wtc4/QEJKqN0n622IYUGM6QCFvXNktLE
xlYk0oj3HXNHbVsiaykWjOqNRakngFm6rR7TLNmhet/YrfqT5tvG7CCrgrI8uHy9y3ZZJOLAjzCh
KdN3aSKGireQSJ6GT69AEuBdoVBjn+/6Kqqg8Cn+mfWr7Lp89oQYtFCVfxhqfZy9045/aX4WPea5
6NND4dlYIYfW4gOnDZJQpa5dfpGy2qGuMqZwQAWwBB/iSt03qeACc6OPNybflqcWgzd2ru+TI9H5
oqHAjcueac4EFSaD1zXBI4EpClSl7PFi6imLMVKjM3qC5/i2eeD62+Q7fElBZppJY6kUy0wRXVtv
zcy3YhoiDoP67QXMphAaRQ2wxLojrbwO1h6vXM2zTWDjg+YukJslrfNvQevQDcUXGCVW/RBA30cm
bGM/JDavU3qKK8uNJDWcrOjiSv8jWSC4vPRNIgmUrA25ltHSiW02Xgs/mE2SBSg9xbJbSJP+jDqk
01brntQziuwr6jDH79MN04y0GQeaXKI+LqhnLE7RPtmfU6j4Pzv0tnZUK3q8a4vqLKIHnej6WE4z
7QuGtJFGMUL8IPLQuE2oRQIaowmCYE874kJdF0zYIhRTGU+3UlG4cGC49HvVfDfAfmx7Ok+DDYZN
tPMMXFmRwPyi5/cOaqFx3MSY+a8eHe0ltz86etLMS8IulwbtqiGE8/uQ7e7U3suiTJoD66k2SsER
FSZvGC79hTIn9oe5cCOSfWhQ7/5Ueh3KMVctwsY5Uljec7zdRkwU8vLm6ACmG3ivC8vpYJXUqdDJ
/ZaSUkp+4qKyXixc5NzlsKJxXB+vdxbzG2w+vdWPuyVqxib4hxnl74lbWn+P5JCZYseImollK6+8
ZKrKZCqcO9pITiuJPNABSEXgogmL1F/Wyuhuku884n/ZoekHAniYhKZYo/hs8U2E95xtSZGxD49I
ulgrGEIQOjvy02I/C29KGvid1xhQ3+GjAIbINfdnxbn0UMO+4HTGuAjOORIaLrRq0lBOF+YdMKnk
YYaG59oQYcOCFSwjmoEkJ9FM5nT7CE1WFOggo0uawfDo3fw3qsif6YmOVOwdEjfEtWqzo+CGvDac
x6hzTtCE9R8lqAsf4X3+AW8XTIcBFe+myvfmofTL363WOWsSVhsOqu0sU8/1KTJcZXik81PxYMJR
0w241LHe2c5SZvdCvnzzDrs7bj2RJp1khVibyh9Lyqb0bi0YcSdirrBKjEawey4r4P0bbQ3jVi0m
rN5EpKYpIZV+weNX5sKO4qOSXS7a2brW5QUznYdCszOh/qSF/cZgiensH4mn5BSXHtXHXFaRaLK4
RPQlIYvrx5Z/gRUptilRiOm1P73qSr6A2aYQA41py+WsJ8grltJAd2Eaa6tAhiYmrW8mmvTmA93L
i0uuYgJLCis1T527mhzycWJZAV6xs8X8mRIXpTIe88AQMNsLtnOv8/A9x+x0pu61jH0HI70ugiX+
TKgWKuTlRobmVlxmjjdO0+jwfLF7hRscvZOFKx00VgbyuCxVjCy3dR+Zmcq2ZF0sxubftMmQ8+BM
W1OXRu5DNmESfkMD6KPz/+aDgQ78gFLQHg16i8UiuaX6XNoB1Cwr0sIpzBxXmj6q6IOquKMXknCQ
eZkR2U0eRgzDXD6Wuz8ZBWJ/iRCf6Kv/Vh6prwIGCBgc0oh2P7IW6eYbT/5vGYw2Zp5xiKItJhw+
pq2PdcYmadlLjLxBWjCKN4z9tbC7TyIUo3KYD6ZN+RXUnQw/kDbeZBlPVwQWaZ411BBTJRcRiIZY
DazyzavPHN0qdYV7Io9NtCHlMI3vcxz0nXmudj5YVetvyMX+v1BJQQjpc2z5Vp/QHwjyDxrePkI6
bS/QDtDuL3j95R0TXjNgcHt+rUjDOdhr+rFK816V6Ojs0J5SDK1Se85jEocyEh6y6l6tHnfrCsfz
buNQs9dTweQzz5Kd+12yszkf6ndLEKNa++YQcTYB/JHVO+t/qag0DDG9JiLHpKeZaBnLEW2Fw0Lt
JZ33FNU9z73e0Efc3IIVBW4fcTczTPHpz890VJIEt9G0pR8DhUmtKG6x059xqEGTudjAoOOCPafy
eZiTUcmrlkXiArnSs0pYAqY8rQFOueicETOlySIOM7G5N+BZkuq5OF8dxbJZXaOKcgGxD7H2CHAL
P7xslY3B95yQDfLiuEoZhRmPFXs31gXls881DOzHmCKXaK+UD0O0RHjvfD4tK6L2F1N12L+8PKqd
82NAxdbjnwxbjRbAJITShrxjjN9eZxjgHhcnFgYr55xxSvLk9GQlduwksLdttXE7Cx0tqpJGKQoJ
7cjpCLC/OamG9GQ9PqQdDq5qzTyoP4U0ErSxnDYknxh0CWMk8r0p43+zeVLIXRCCsu1gD1ghYMpR
JG30sKWi1pLGTNqsVfxgRXgD+h5e3jGxyFZRSS/a88GeprNFciws/SzkDgpmdr6m1vhTiGRDhn3k
PD4Snz6hCqV/k2nwNfOeup1WbXSN7xeqzasoV69Zs2g7W1/zfCVKfCDad8bXKTJZ/GK01EhHe67o
Q3EMxaTKJ7a+lyiQqxSz12Xbm41SG/Ja4mdw09W9BZdDSEu6JQwDdPojcg5sj4c3oYKiFJsnkV+x
4ufgkgxWa7e137dLIYLPmkXsPGIu4wruojO7caUg6OFFEIgN+17AklpIZgpE/AZDMRtkP+ZlBqY0
xY2pS/rIqSKQ/CfndaFP2i1sJqkGtYVDiOtkXvckWJ8FBd9Ou1BQYeQBjzSbI6BzQymFvdhUkjtG
VAfqPgeM8M4xX/sWL6XB4CjhtXucCdtiph2FMKuPFdjN5zQt/poZEfF1nugTOaOj+PCAbXHvHsun
ifuCx9wEi3daQVpjf2+6R42eRWm5tVSeMFLkoZODXKXvjEgd/9ViAYcjSqYiWe74XGXfDF3/zzn4
tV1kN6yC3ddikYFBWoTtGn9Fpbeom0KUy3aqJ7O/hEUbzB67V3q+wi4e8PC8CoPrUdWeNoB0wIrv
hP8Z4QezfB8ClCwVeyM/Da8SMZskoDT9Ubx7yXt6PA6wZQAjmBFoN0TcO3u5lC4pdjBZaDcRIlLs
dJNk5zKf1jaTYL8YyozJdGHszAIIRYQ9plk49OJALpnJ6L1syUtsPpAlfgMnaD/hNoPTG2T02BwW
EwbYTrZqtChye1/6xvdDTwsl33ZyI+zEIWirHnPNr1CkWedKuGlFlx3T1/4DL4eXf14N1VyBJawF
B4EuE629MtBf0GzG8q15fj7WGyEckvylP/tkXqsvWAd0UPCGxLa6wVKCOhugmPPHB4W3YnFwBehp
/Y8QqiUeCpnPfAPabH/nfh2KgUv8+IsOz4Na73sOii5fdGG94H88kHlRoTx4PFSSSvTBCThj6hzb
kOOGH9l/XqIzsb/hAZJMLjiZiJs3u+VejpBYJIPbjq3YICaS5ETDYmTaANfDIAva//AfQs6SqloP
vA5qJHLWVt8IVTita7Mjv19NfBAP/7HHsTvpVfKGYlAU1NjoQEkyKTJwFCWWML7C7R6vd9m9bEoD
Eog4yMrph0qnjfbw0/qHnl6rwlBPB1bwoIMMkI2bgnXViO2Cg+XG1mOZDziTai2iAnb0dqgCnyar
BVYMVqWh9MFYMijfD3k8PmHDxviqX2SJiw64YWHn+TGR3QLWV2Esf9ODSUbDEmtvv1tU3BcBFIZ+
8UT9PO3TW1HYpCMRAMMB2B/KlzO60XdYqmU19wUhW3BvhMPNu/i6E37HxK+wCrjOpnvjMsWwHtqX
dI845tIQYi+0+GObmAjtE78/S2iBlZT8aLaIY3o9Dq4aJEKqQXWC1IzqXM5Vl+w/PCwGd7wg4N6u
wgJ1q1iN1ejKaGB18d1nvQwOxHpH/gjKUNyJpT+g7OW7YPxFMO8+37McSud7RDZ5VQNMJQveVb96
CpcBPb7/osR5AtAD9I3ijzCmHGHSKRUDiH2I8ETEVsmhysa3pt8/0+rXhv/800Nu6bw2ZDoZHXSh
HXDX30TTRlN3pjOgaIm5LKWwGvGhIT7bFR//Pr9Im/bTL0+eMramI/frmUJngS3s6ue2uyz6/0rT
H1CzNbIevu05igIHEgTjMfKmFf69T63EyvYVXRWluXt6Cdq561FYclvH66yE9sHMDvAeSEV1IyWn
16B3o2pVhJHlf1cS5WZAlvLgOR8PJL9EgFQCmvcfYBtGNfVlPCVyp+ZeyBV7Ct5Jr92g95kSbtI9
n9T1TeD2+0K8Ym4+sKG4qvd7yCOvmx2avDKAr1O1l19dYoWFwvC5+EL1D+N8nzCUSPy7Ti877WhP
FGYFoy4266noWP1uC9ASQqDyEERTFDBrV39EDkepMyZ71DFlQ7eKzDAtf6zdXTQao76RgVzEuqpr
WF9kjhDPbLNrP1QTMhLgZfXO+ifaG2uyTYJfHmXkaLEZwTnXPq5A8Y21swE3kuFkszGKmzWMjlub
VNPNueAchK1rtqrKQzJ5/U7OY6FpOpyuyaCxHvcpuIpbsYaELQW40nkiIlMMSIA9ppEhyRWasog7
ttHUYyX3MtooGB8aJKs6lFEIusqhrjBwghq55GtWsDYj/D1ewTRpa3AYK51b4C4AlL/nBgs76Rjy
nN3JSRO3YG+5GTmuPMDZNbAIwkJDveI0Hi7cGDOujQBHy1nFfzNlgPu6Owu8APVcYMssXKtK6VAB
7ohmvNZK7sHA62iIfzsOd1YcRwwmrismfycC/RbvW77frf0lxIWVLqC6SxrRjdYq6AZmUF11ypPJ
i5Sumn72VXw8e47Ht9suL8oecfHgji/HPy1J+Z4bFB0VuERiVah9d8ipVz8qTJRDgIPRGxJcKY1c
da94IBkbzYnPtlG03rFArZ1ebDC9biK55kapYHDu/HnLeL2ZNzcNSCfTj1UZtOIJIMoYp2W1MiVD
wB0RMZdQqyu1QjImV7bznVX+iJHfjkvm/fqZNPKabqTwIMz0uOKiyCSgVYdVI/+j+jV7lvGmB/L7
uGAwHIOpnRQh6uY13jjFzq41dV/fVUJ8Ct5I/TZASk6itwX3qfY0t4+spOyuu731qcxO47OUS/m+
U9jisRsu+PH7Xjr98vKg7h874eoMxaALA9vM/9LivDN6aSmfYBc8iBJhE1l1IO+jPDGNmy0mOIYj
0iVjIB2euxAZ0ZX6I3ESbYqBdpRcZnddSWA+ctArl+viGBzZ4mQyaRYlobsSX+K0bUaEBy/lhhbD
xqhrw8G2BRO23A71m1hemXlBBc+0YTIN1d7a6HUH91MQMHFFI67uf4sN2NleqNtPPa3zlzFbeHFd
FU30qZEuDmYfIhjimXklw2Sa+uKx5WJdjtK1vzMNK5/mg+Vtg4TSvk87OhwBuAtTTjbLdx2pklS7
YmppuqruLrMY4JpNmo7oTzwoUZhknWrWKoaikLysuGUKRSkc6CXOYCR18FTdOUu7w1CvtsJUB4BX
FpwOoSHyBVEbbnFzNlltHE5BlETttuOOrhN9NyUXrc8ucmE1A/ZjOD+mavK3/zV+UuV7voJm7KAY
NZnx9aDVsvxGx56SPvaXN7gnDFAO7DHSWqj4phA1m6eiCTtMJh7TjTj0BeCBSgaL4wMqfLSVf3ML
pqGlhAHj6qdSndgK60mBhPZXmmH++dChJgb6j+/18cjisCXH5LyI3+oo4uGj3Ifp7om3kFavsbX3
cTLTT0GJuGxVRZOV6URdtvV4nqmjbhwSc4LYIy1depr8QwGL8Bq0Wl/dHdMCX/mR9anqUFJBeiu8
OHQZwg153u8WDCWY/ynQ3GWkeOAOwv2bPLdQm4i25W5geIN2dm0oOeHcpXHFVWz62UAyhSaobsVX
q0osLfUWN9VURmwmYEWIjjJKueTcSvWiYrVOrUdbAE8vec5WsfmHNvHd/09kI7Utid8evq/MSWoS
T46edNPsOeidg9Ex2j8Kz+Uzilf/7s2GiOZ6ZZuvIdEj/TLPrTX9VTnwsvmZ5Npjfdvtty/Qgnd7
HnxIEp5c+fLu/UQtmSlkn+iCuYyyVSyRa+hMoKUciQ6J6tZtMxVV0+4OXT6kD9+d5lf19OaFU1td
KwQ3YnT/NvZ7JErI1O6lxNlcM1OFuu3DuxRLQBxHTZq9ZE2VYiCLwFmZj0n6COrIjfT8T6WHul/L
7Q+lHQQ14I+prEeN+zo7MozqJ5syBbZ8GUxlnBXS6mv96Ek1APJj319N1+VAA+DDH7BEJXLa/2mB
93MrL4IlFlEComyy9ctUG+s15ZVgnxUSGQDUWi3KXL0i0EqTdFVWsCn1Gynk32L1pCzMY4bBJoPo
pEFzhBSmGM5ubCrgFfQaaewmZVNCGsfl01axBL2ftc6mtTga9sMgvr5496eaKQbrfMFWgI1gATJC
Wv1dhexAXHNplNyJZzie+npBrg+2Ool114IeYVPvzWPJfWmn4cM1ltWGIcm25LK2reUqIyvZ3U/4
Yzgbx1r8FbEIZlCDMsnCO3wsInPmZhzueENwzSIPATX4hZfZ+mBNUBXD2XW927nJqO+Y74AVcEw9
Lto7YanbPv5mHFfl6QWLm+N5/75wd36n0+7+0cIjAQp5z3Am+iUshXbeG+q+Pk+8nrea4u3gVaBT
yZ2vnwiPhcNvaMnjPXMWGl/umMB3T+jqkqnBeqfiAuGOkRgqq6JFn2W9nWlKf6yWDij3gx7u62ol
ady6i3kTNErhYevKA8RA2dnvV/MXPr+5oummgzxYN1f/vsLnZqclmIFviTBh0VWJZGhRvC2hN3N+
z3hq3pkCHOromrZYLxkWZ4ptwhrJBndNHHG50R40UBY+94OUJmr2Fs1whDnq/eTkB70RlT/PKtvV
u/3SUy/bHXImF0m4CuBTsyA/tr1TamL3cUFPMtPz+tWpm/mrRxUze1MPY3uYVg/xrv2NoaF290Y1
/LrvGv5dV3tekfmq7bTcBUNZsfpxxozk67u4k3O+hQrScGR0JTFLlU6Sy7f7OmBsoN77e1iEolmH
zNEq8IyPjHhW+ZQlrHJ2zAe7tiajG5N0CGPcVw++9UKhxj6oOKFWisTPqm8TIqRh8mdRAKOcm3tS
PFPS9DJaPUowZUbCEc2RaIAB0OF+2kBYaJ86tyf0yxgzvP4d8EiBXIQDTKNaYXi1g5X2nUK76b3C
WHL0h/kW813UMkqsH3tk9sdrSYVi6fKjdrjx63kxDi5Jou+Sg3h3Ovw7//YkEzuff0Ex+8zBIB/q
w4V9pc4v3zdr3MVDU7IEvyhDrFXMt5M7qCQujS/LfMI41SYxrlh0yjS8pl+r+pDOyl3V5UbouU9x
3yPYtC+3JiWSW/is84+VtsJj4DI/5/9n3xPrLosy45knOGt6AiIgImBQBpdwlp6spn2PpKONZVm5
0JNCDA0MMrfqrh43siTewAqbpIf7wuGEACLG/pmu7ZECt3mSYYpThX2h8jfCRwukD/0T2WAbQ0Ph
Wbicl2YU6YUyrr1dT09gZveuVewQIqpP6HFJiXgkrmK/ltI3vpKoSB5ht8I+MAHY0WKMmg3eF+0H
ESz1pi0VCHRmRdbrYsb0GNizBedYNkJTntWHWGfjgdWi2bONd2Ok54b4KDp8+cZHRfSVmgLnC/5j
KnqhaFj7GruA9nvD2o3VSl8Cv//1MLy0gUTUE11o0y8BCDvRYpx3nTSaLaknNVka4c6jOv4j3kxl
ajvSSzpg1dvTLi49SAr6BLkuum3k/Ej00N5F49vHOKOU7kzOE3shT0gAATO9W+gJgaX8Wm2kI1mA
UBHSV3zaH473CEQ1retiHDcGTosV5KKHbo5oc6kRdmwTsV0sVwbqo/+ybbsLPIvtJ6rZPDqKYj9d
C7Y6qHvlzv46WC0aDfcUuw2TrWZYDFYYCiEwjgpfiHCtQFo+7yeAD2JfcYalSCCfwf/g+PbbvMXK
2UHvsJ6e8NRvnkt6bGVZcwGJdDa9iVB5T8ZIOcGcs/g9MpzmQT12FdsFCE0EA8y1MyevFe+GK83T
gZNNdDFGq76lFbjKrcd7dEk3mMW/pRSi8dwYke2wrE4pbQndZ+UuIWk+lXDgfDxmpOHA9ekF/9Ph
tWqDGtonk3tLzUwPdl2EDMwntjZw/yCm93aAZCoaap/KFCmJQimoDek+FGroziXsumjxcFnDLoCs
EifR5fNxEOgI/0E0IiAFieGC1regrSsWsX9soHzR+toDksVIofAeVyGzOtRvCLXQtF/NagyiE33/
Uo6hBZkP+Vz6+SZCiL8Jl/W+SDPiZ3ZDktx5rqBUMfr8GyRJORiiEkjcrVmFSOMH703x7gyAXNdq
OKRvHlQoyO7Ci7sJtNkLbPnn/dhGHevp9XtUDj7RGMnTRgwdYBjPD+i3kIsfFUhSo9tl4geIuKtM
ojZxMbAApqn4lqtP4cObdlZvd6xF9A31lNovfplBosSyAS6Z+LeCqbk4GkkVsgJ7KjkEoOOuxWch
f8WTBBeqk4atm9HJ4KtOH8a8LWrnV8L4GzGw6sjqdJYRFQrhRjxrE0lEkxfBM80RaFAVHCeSChRO
pq7tI3y9QhNO/grEhOi2AP85Bt67Eb/4tRcl/S67bqxwlzZqG8m5kPWWWQ/Jl716VISdjlMmFOp+
87aJ3fhRlzDyKPQM120dpqWqHJP8N3bgAkkqdvb1jSDDk/q7VRxsbeS0GZ0bAtr63AKEZRI2xhSN
wBIN9gwhogp8Z6CZFowEgFhcqEIUXTaCpCSnIdNhUVyfQsduXvw20fZCm5xCo/4tBvAnVxfmzRBX
u/4L6bPO8A1r2m2QJlmuwtjeAOySj1QN9gdx2+P39pKnoIsnAI+dYv4TeUfnmBrtU6ZUa21sKz4v
QnTon9au30Q7vK/zqp9CN4Ajzvgh39XQnqWFcyQBUCduEet9qv/xvLbjEiQLMwk4958Q3ajbBy9l
uuHYr2dlSoWMIoDte22Es948VRGk9R5sj1CzuEtCDA86tZzkNuItCuSX7DtzGWHNgclE3YYhnsuy
4wSUhhShOZbAR7Q9+Gnof2/W2OM5gzd5mvQEERwByhW39i2TaDHMi7k5nXTCc74fa8I97A3YdmaU
QUvgC2NRETwRb6qilHGQisHolNbNstNof57ve9zkwx2PnLHDc2EIZjTm22IvoAGOLW0z/YGRxDsI
k1sCnEj9M3lbYP3Tq9HNtufFcb7iZE+Zo1wK28HUocxHtfcW2M4kiQdZM+fev6CJxCh1T99GhrsG
31QUdFJM29kcX9ycmP9CvuCtXp8OjLXiI7zgzQvqtz21g85RRsXD+4WJ/Uzdy6C74Gol0O5OvzQy
g8OpPOPGKk4iYI4Lzi5Ib2WDuUh3gy093watcChwFfCj40cCVIO+fcKyCIN53L6xR4uO/ZlEp4wM
SEYRR6YNdCRCsolaXF/1dNVQzokLBVa/N6JaVQ3Ty1bou4Q9NxlQOo/luGhs5CciySc2J6x59uE5
LGYf286vN/7HdX7SLizws2MQ6E1QX/mjdejoK81mVTIOryP+lYPjccfimjHH5xH796OOJIt0W0fJ
t24oC5NMQktFj+J0unI9QSc+FwbORjcW9Jkutijdz9ALbW/ISJ6Oc02XfdqajZvu9oft2W6MtxeL
icN/UB9aLA9geTs+pCe7EAv1uGyIgURI8iCQizb3M6lHgSx0sc1NazZlNP70+iOEueDWBgpxhH2B
mjpsmQg3vPkSv0eD3eFYZxcDJfKZdFaC++UA1XNj43TVsvNz7bmfhqQ65MPbrVbh4EoZ2KGY72X+
8EO8wRURvUejkgKjo2a3sHsHCEBYgIsHpIkDb9EYy5pacfWBe6TGYIJhkx+GsW9ychEEWVYtpjSN
ZJCioBrTlK2wq5k878iJj7cjH8c82t/Sh37VpimMkopTjvC6jA3HyCtzulzDGMietu6RVEmiMpzp
8di2Om+4Svtt2A7+0E69JteOVMJM/Yazs7R9I+uliUs1deXh9LLgQGagWzxuMnBNcu+Pq9Ec9MPG
uZNKPfqUlDj4u1lPAjg+54pJp8x1hR/Pw5e4RVegBT7WDAYhLkKnrc4OoqqPeqPpy8aOul4RQzND
eYw+efrn7mVJKxdBSjfORUfc3kWwN1AS0ahN3fB8Gl6psTJMppLGUL/+0RovDkaJYPJGZ5s5qOw0
96pX5IvE8Q6iuUMs0P1rFI4fDEpZoJsSGD7RrPsWri4u80El3GLJ+9nvRq7Io6LzFn678m16HyKw
O64uZG6BrioQiL76FN3Vr15WwU0M9Pq7LRmuMIbMFIUQXvJwmKjFHcin7gif7cAkbZOoyFOXi9G6
4n4kqP0Ebu4V0Ev9v24hZ0Mbp6duiOyBS4KM3txmtP/t85nKXBsyTHhPoubdT66EGPmqdS5JEhEI
A98t0N+aNpt59pYHZ8z041Hdo70Y+chnzvaEX/+r2odLvCzkBefUoiUqjP4nVEvZz0Lss50Q9VCV
0ldoULBxbBC2ofLVyuHQokXJTfx6uB+g9YQjWTF8HSPnKzXDbQlYc7X9DeHDiOt88PVOGZC0IGIr
YmKffgSVqkja//lfE8rh6BuR/wnLSR+aU+r4ZkmQz5zC+wF6oyN4TnBQ948R7boT2zikMIqnA5WF
U7zIGDWsn+NWSX40VUf3P07iJxava7+RZlhByj/5OAb+dbGFw3onExYNROQSa2L8VvBjX27BrCq4
i5kRL71ZMTbCfHDT4X8pMcpkcUO+iR9noyLOaJ5+kGR9hfNXqyuoZcjeahBI8bFC1UIX9c7wMoDa
DNqkIphN63dELtCJ9arNnlSBwL7Y7MErnF1jgJH8Knv512tx1ZgiqFre6IkVBbF38DydoKcemD9M
Z8SBli8OaoTXC2fghmMqblAaez/yB4f/yJCMtzN7wHydWY7p9e2j8p33gEnm2lciR8CjmBOAmInf
pYs63i5JvpT0FpkfXdL4MCVygAoXGPz2IRnpN8fIbCjB1+Fc/q8l+3sdlkyaO+q25gk7bye6he4K
r/tgxo71m3GBqfLlujmMrZxF4JJivCdJZsWXyyAEc0xW8nmqidIfRCYyLV9JgisPZd/TZkxaFp5e
SYmNqZ690pn2HwRR8SR80c4XzI68GT9uFVSacC5EGBRYFTKYOnc9CvB88R+bqBnBhdXQ96O+F7Q0
xlK4Kj1pl+3iOEbTws+LSO3dIdZba2VoLiSNCAgCuV/FoXsAsA8qBXv0oBd5rI16C6aHxXOZDGsh
M72ArsvlEgs2aOTmUTXzM86jHqoU4gTc9Ume0L194FPsXXbXHYX1AGDfIExNiVkDXsGWgyKoyRuY
974LoGpzohqcVk5zaHeAP0ZiW4EVUJSQKBCDq5rB8t/sZbK6iEYgt0aH1n8syYz6WOUb1AdwQkaJ
ltVYoy28+2kl/XRaUUNI7QA2VRXEyhDqNFZDhBdOUele1HVom8p9wl/HSChiJN2EiqkaED9CapxD
8uV1Hyv+ot+pp1G7CU39c64kbLRQgq8rNapYWrokHF7vkbV9WB9ULW3zX3W8ufXP3/AwgGaGUwnH
TWtya84DnvJMbUzwx5Yygi492sEDqUlzhdSFMFvJpS11/btJmMB/qxs1FqRswVJWlM6Q7XNHxyMo
TsLXzGn14up9X3kwMTt/ano4xzmDOlMkSDZZ2ubacvPsOKt8cr19WnLuQeBnirSGadZVnJHdaQC4
HddqBMFc9K19EMUjqwFlX9ikh6ECXXQ9E5RpBD2rGqKU/4SOby+60WfQYO2CAFK2r1tJUUgCvQVL
mcUn9guAPf0VRMHOZU+46KxvykomRBlGSc1Ol6txv4VQnrguyHX+U/Vc57h8O5QSD5mT3RIHgDDr
ez3rUalJATt+JC8zl15+Wp17LnE7lJjk+kW0+cuY7WteUrhRtJO1tWo7S1lXRLCraodtL9OTjspU
X5+wBa5531Swlo7CMsotae/qc4hQH4zzl8taJWNLjd4dYNJvwxJARZQJcQOupGUi4jxrUWgNY+Hg
+cqvJgIjRjKXU+/wt5D8d6ZKAmS4cNd7tUpHEF2stZc6IcAaf+4wcUVelGPbvs5yTMCDmCAdNZaf
aZfCleDneUGnwyiufznJSJoBiEiKD9O6GMrRFCzBl2bjKuyV5GdWpK78g7aRPrMYgouH8k91uTld
WUzRKbCsr7zH9/lvmYWV6zcOBpDo3TNXVzDW8V2DMti3vPHbj4MyUvgBVO8Chz2XmLupUhGCMLY0
BsvGCF/LVm1dkWYN06DPJTPvAqENeoohSxwdnmRwOeg4gHaRuysx9ZjpSzGEHfYp7SDZ+0qQE7Zm
u6ZHSqv8IQFIBmYJhx8ghsBR1JA7MDxtOrZUPl0UmG0lEbdGsaSLLu9/nYjOO91wrk4UFgxD+6Xj
QPeRYrS5AjNkIMwJPiKKTcVcz+zTYL1pp1qtni+nlEk3WRTcjkY6r4qnhu6tvY/aCojQRvEZ59s+
r8Jk3Tob1mdzwUj5N4UOB5KHQcv9lWdfiw5qb2gBC4s3gtzU1R7I7S9kZjx48tUDdB9jiTv2TM0o
btveg7mHmAepM5tNZ0LQpvkJRcqDwCfz1VxdVAVQQdlBf7OpYRw1TgZED3me8CoW3/4X9DnE0YId
/iBXUS1Rd3gfYIVb8estvFjNiLGSMYjvAOcluIwxggRr+Cg+JpByO35m87OkgcJKNjSmLyyb2q3r
6zauJN+LeswPmLh66fqiwbcok24SinthCIW4v67dpuUD82k42BiysqNYP2S8T8TWXacRJnpe+vj5
aJlUod9HLEtHb73B4gXxZU75aCDYHqCKLrAgJQVp77ZDe6LaFNSHENSChF5v2VUfrbjdYMJh5r70
G1a7yFuQ/+BqsLDozOcfsd2UJ0qk160gp+rbyml0mXe9gOvbc/VdMfjsReU99zV/zvHCOVgGmSxO
vZhzOalVg9gHFvWlycIyGdnkb4uOFmMg0LgeGzmHb4ZJfzxy6NvCdoRGu9mGiMS272i5VguQkRW0
IfQJL6sK4HNiI3Xe0U5YnjGUrQGxzWqthPET+EEJxTVmmaL6z60zIStrDma4+M2Ts5gZE2lOu2H6
ajIbcqaAQFdJlK6c7hBEtWHFDiDKiGO2iJZGwLI9o0y2L+/nvGyAy4gDmBGCVXnMnjwx0hPwS3Hm
/1blJbEW1mxowvl99JJ2pSVw097TlKZJiN+yPsh6PpSoGxnO5XviQK8SMuNG5bpf28iw0JXHbhvX
w1OZRVk0OCZjVvlSXg7ytPhXUMiBDlzsckc+wuaMj0MbQugPThHoFkUGjLlls4NwkWeVmTAf8DPa
BJreMi1vH9mjD2PvsWknvm2lN0z6ncQi03eWAN0uSpBSZObWv3Nngnfm7FVR+vCRGYLN+6e2S4af
H9SFubq7seDnyEbDRq+Y6ITWL1SglgdvtyrfwNKtD5hoDakE/zO4s41hAi0bWBxEc3v5HQ+6sr1O
sc+hiCRRPVu1ajWlKm4YJ+QLoPFw42w14ZpXU88UAcRvKm4zKKPz1MJ6muAri8Mi10SDmQcMF4YY
gVUBLMRdk7a7ZSwu6DXVO6HZpT69zjSGlM1z+M+WuNqWavbTR4RJw88U1zu6m6vnox4ddBOVDRM4
oC4EyVpmiLY6ochLLOFIbkXc0SIn/qReawh4P44DDnXSCU5ME0EWuE8uOpbezpdzjPOcj/uQx2Oj
Kmzex4L0oNy4Zv9COMuBum1ZxkyJGus6wTQXoBcUqVS9WMUDsOnK8/9VhpzlWgxVsL3Go2BXrAOi
90CGmbxZ9NH5/tQ3hviFcizFa70N+1UEBiPaThOr9Z0kYBVf/KhbCCdQJw05DEk9nH7QxW5eMDEo
XBqXlvW1eweK48Lrco4v1+p2kjSm5QGlYiguH2+F4t5ZTkgnY2Y2tEZj2cJlab0dIyZ4U2RI7A19
4zURpnhL56DUivY1PYX2znE1N51uanuJiEJgvTcVmwYgXtJxWDyNGgOxIj+fZ9vnDnflRL/gPHMg
h3xaNVSxsnPuJ5OSOyk/b/X64gnsntxw8jQPL4Zb3BAx+4FSSLKrz/GGXbGpkRp784TLQXEiNCwg
nqxMN+eCUz53ZtCdXcdYAe+JBdtkTqi3DPiClZKTXu9CgVMiEBiRT60geWE4zup1h2Kp0TXlvonp
9cet6YifSyOJ/Pp2eAbfciumubnp3Whs/HPIO20W6Zq19hWklKb0okUYWnJ3VIXbuwzpMN5AZrIK
3IpUxh6QSOkKf144E6i/56XzHAkMH82fRLguEBm3HnntBAHZrJ03cQuxAxSo0dec0Z4sbjXv8YjE
rivoLN6LD7bHtcm0o2hbLma+sWhtkHvBZUt6pigc1UD5sKxBMJacEPE6Dp6wccphue1CcqJIzaM7
1FR5sVC6a4zmZCSopom1k8gaAtnyb8epxVD9ueE9ud/dZuTG/wxH/N1ghwaBKn9If8bvrDUrXN+B
9FYo4clQ4jNlmd+RyIoXPMQrYGXs84wRxNZMUynOI534OP8DRQRqm2ZE2rnc60uDbnb0OlXolTeO
2EgmZmyIQLju0kIiPoDKeAiXtXVPmGhhfCra7UXRZCBsOr9MKZSJ5C3f5MJta3nONZUUH48XGGtU
M9rsD3egJqbnWGxRxpai9KDaMZT2zNKnHT9QOnIpd5NcCzduXL2GZ+XCF3vrISctD/8yeML+kLhT
pwDfzneFUqEavRDeqrcjXesWnTdUzIdo/JXx4+SOgYU7BNBFZpgg8E/JmqH0WzVwcFRb18YxcrEe
VJM/6ljxOV/jliOtdYQLvHpAs/bDiLmxwThsutkqrL30ZCyrjz/9vm83x7y1d7SMzlHCALjB053g
PBTsbvhasE6p9NI+V+l7EF/WRoUZd7qm5u2ec7iAP034bY1hAeabOYru4/6ej+gcxLubUyltpijg
ABDy6H7/SnPY3D9zqA7ac0alw791E4Aplf9ac+wm8LXtPHWB9v7j6+qD9LugXUwHQM1nvaGjnQM/
szEllHDw7qrjKF2F/gdLG3ZrSbTfOcglenAIsBB6PSv16NeSsWY9MaGAMBepfe9fiGpDxANvwPa+
YVpaBnzzEKos2x1qFsR6K0xsbe9gjVhhZYsGOZbUIkoq+c/P7KxDlGBSzwZVi+XldUjyUvCOuPA6
DgrK2ccKh3LnqU6N1a6cjArD4TlNiLbAvaLYAwqHZB1CZLoyoSSZ1H4GUOceP4iEDMqpqgkD478+
odVX+C9UQ3qVM7+ja4bHcGjoQGEp8XWwpE7oZCGjn6QDyehztaQer/WUd0rfejzg+hEe3sCYk4+d
Z7w0cVviGrB4OtF5cVklS65XyHbIq6HT1M71tPySvuGhtpg0bzE9iOp924xHRQZpYgelZpGlFnYM
GmG+wB+/x27Ede878gIUJMY102EN0eOKZhucvRzqmD+rx5gj7cmBK+MR0LM/o0f+Zt1gdqnBoHni
4L+3Ba54WtHvMohVNRI6Bv4PoDQMT8WX3vKDNfAvkEaH1ffV5re/uvKxlzRqwBh1AVCEkX7zRyFW
5w9yxtwNaIzEnRXuKY1/rUpM0+KzIkP4mpbL0LV2r5vV/8AEhVZo2EHrDjJf7eoIbLrSeWdeQd1U
2/ePNSSbDbRR4PQC74vm1kpizcDOm/SKUMt7OzQ69ZOHsROYzGi6QSIN1LV3oOe/5nFfIWyOA9cP
QwaInoAuDfjGMfwE78VuhB7+nXXeXveGhMVM5kC7VfZ6wX/rdsIG20cMMOkuhmnEWkkKdHxZg46w
y/BZKz2ZsFwBn/9tjD2u4r3a1OJ5zemwn/O/f5SfusvxoOZrjhB3nuM6aHdJ9H4W7Ao9+eoOM+Ih
8uizXy+YkHz9BdDqTDp7taQXApxFbmm3qR9qofprdd69rZPIobwg8PmfO/DUsV+VRhnyn5nMLJ15
gSNaPUf7FnIa+OtTx3Tc2IRDLY8K8AfRfOeFTWBXVifNl/dgh4oGK6FTYFTDfJibF5fxrkKXtUVK
L4E59ukekq2ulbqTdz+Ri5KBFYa2AgqqoeEfQzR+G8s+Ysr3EU0y8teoZSQ2jVvp1Jwk2RrBBfoB
XWt8UO1Ghz8lcwrXipTAZxgkzfPvnb0J1HDb00d5j8v7SpXL4W5xt4qcqZhuph1mrZxrbnfdI9uX
n1IPLIxl7CssqHF7KcpQ/htKBk19xE6DnONue42ex3Q5cbcgi3DzbQbMqoiBoLOvhyzZ5aiFAfCB
9VGCXJuKiF6tV9N8atYZzzuA049l9d83v6kcfAFmsmhFsVRBoO8Zs3IwJLQJUks+Xk5Vvh/MsgAR
IV2aR1JZjoxI3dtB5I3K77VLS7fe/Vr3FpDCYWuJQ5WDUQF7B+3reu20Pi/CaHw6d0GNHpLh3iVy
TZ1CXm//PvzTAjeC19UhvznUFbKrlPMNXif791l/gUDr4Sj8Vi/STkMY1qXoY+DGcndU/hpvZnK4
Ox5FROYqmMMUL/dtS+Pr7HYN4WsY9TRlOMowsokJaoM6OdO3A+np7E16iEkltnMvwBWxuk8A4Rqa
pikzncBv3LWYC3yQEEq2+7Odt/Zn4WzH2d5CxISgCpJ/tSwXPhJiJFPQY7O/Naqmd3L3/kE5RhlK
WzjU1YgoPcvqFiAtsmxKNwNOQJdB6Vyvj1k4rGw8FJxRlglhGrAG2C4Bi0on6yAyHVaNG0PDjqNZ
yaQi7Jtip0lG+bvkogcM+IhoHEbhIh9FNUXnj2f6MH7A/sn5+Yv6yg0ql2WUoQegE7tka/MXFZFS
HVdExxKxcN5I/Y6JF/MWJKAnBaJsH7edYa4NOHd1nPbzzADfKvjU+0SiXhmZYiyJEKhlyBYl2yll
SP+nWqm5vpyq/ftKMf/dvq/NsYsrvS9kgM/KGG0DbrQbHHaCsCg4L4HNOBOGlcThWJPGpaP5nt71
/JecOXu3BRpbZyG3wEZqQ5L3u5Vsusi2R/7YQtDl8WKSMwbRFHJz93Vfym3+QsxM4A+guTPFBQB9
jabZIl0Xe/pFYij+Y4HHtI5YOpBdjwLVVw7P6lvbma8LGd7/OkxcOlqU9ZhMfikEvLBIF9aOxaXx
pbFUkruSc3m/kpwfYxD5e0pXUwlU1tBFjr9/sHwX9ubcOd+K0EYqAaeJcD5Eb6aEsEMt+ANLifAy
E2auumiEZlWxhwUPuhbaDg/+WMTTB2rDL/MTL3gTSnthvXYnHpYW3vJGFpRLtMFzDAh4UWGHc8zY
kDkFL+JHFW5Ihsz107BghqO4VZGJyLAcg4vHvUfm/19/L8T1diQx+ei2XvFVxlWqzSjGbW+xzJC5
b31eqk/JjoIMWIKNXlbSFhOyuviqA7QGBPPMPGj+ipgTujCZxq4+Aq911Vfu6znqUb79w21EfE4o
fsAoBCUnhSyzWx0F+cYHompl40PFsBfRZN4kRe5auCkcz3BvzGZ6TDg9XxZ6t301k3noK/GX6VbD
ZYAXBkv5Tkir53HZF6/nIbqOBxFiom0Jk5jcALhUvmt0cs8SBKbD6Zcw+f8Mj078finaGLueIX92
2hQ+BEkndFV2BL6s/FNi2RRE5hGhFOXLLYXkiyURBXLAr/ZAMqdEVjUtmduuwzQ/xjgJesAo3kGX
Bs9onjClQgEXqK/tx0mog3VmGQWP+d9v36edeeVUyYqNWi3o7N20YWddZ0eNe7moczv6TLzFgwWZ
/xyHrrNxy9xH7A2ih/lHAweg8QrLcOoyQ5w/rldw1VHjHrnvfGLs3jyg7dnR1IkZ/NIGp6s3S8qm
FJW9Zd0MZjxXB9rDhmMpr8U86v5aGXIm+yOfLl4tPYDv3ao/4xgKkxPWzDKtvZhq6kFuQ/MRH8gL
b7onO/L07S0g0rEwT3rVxG3uxQV6NEE9xUjqWeM2+1EQp8UV2k8lMP1kaxdt3t2m8CU2SxiCY8P7
LFqy/IXO9ttWoYOoZ3aWMZDMl71vYy9aVGD/fr19TRwck/eUg/C5WkJG+zKtylMQlsIIbZ5iB4xs
dg1ijQZ3XjW4i0yUbl9PPoiep3h95wVKCAjb7PckUbbTauvu9Oy58jdbX9S1hxykbCm6WKp+9tDY
A6bopd7ldjhmPXhgxEmIosnd6Ya5G+Ej+RmSrb6dKAfy0BQe4TjIAGqpV24CGTIl3KEY3Jih9dC7
0AtSPFeZ/vzNGX5Jq8AzvVAy35WtgCzpdQzYRv5tY6DNkZjURk+xWkhJi7R1LUjd+5uoVOud5VQH
e9uBlzmCBCZScrh7sPsxouBelPTlGoJUhnM8B+uWZV9h+4tqHEkLPcdgzbcjuiT1FCrCLXWTUSsZ
2N1W3tRw40gtiqt9j3qW8UprpkGFga0Fi/uritQTeZBTFs/5/qRw1jLAm6uEUVey9yzI7wCSeAV4
dABfxpWwljXLnguyVdmGzDbBluQgCevJSFpCBknAsPJiCXKyjlCiFvzgklztltmLHKwK90laxWuH
Qvlr7Vbhfn7VfWRuATIGiRrN6GVmfykVwWrkzxrQ1cECstrDzHJ//baWT0vBJKA8K+OiTw8OKGrf
452D9RarbreV0xpeUdTlmnf01g90ge+yUSx2hc0vdYM8M2xxwmNMeFaDqO4jVafXopwfCOiMVVkr
0KP0n8iPt44+YtNNM6qrYvaPorwnuShRALgHcsYO1v1p5dGoZhNnU30jh3bHz7qQFK0uu/IkJ+u2
oWMlSv0sDGIBNdjBBCgw6/SMrmEsHz+a+/CD10VYpAP7FlAxwIdEtUERlOAuh/24B3k1hUv1oO7L
yr8eBQ+qnD4ZHgLLlP9QdA+Dxxlnow5Cn0HHxkVT4YahozX6RtgmQohLK7WMZpGiGa1HsZByBTaP
WBUJt/bPYZwEqVuoUBP6bCHuOZ8IIvNFTIb36dtpXDHNr1iPiICjCMkcywB/uH+AJwq+fJUlnemW
AiOwC77upGTHqdt8sAeXyu1AUAl85d/tCweU8BMTASRlcvPFyTqEH9K2fsk7ilDlKjf6Bc5bsGWx
XGPNqKjdYg/2INkgP3SLxZSt7Tbtz0gmV91p4T9gWabuL9OI3q98bwqMemUxqq0dl1Eq3EgDZr0v
P7QdUjRv9Y5Z1FiGCQPCDUj9kEsJG1g/TEQdp0A+6H5WBin7j3kZZm0v+zNwbKYea/qqpNDDXhpB
fUoPotbGzPIY7H225j9W5wwputzACpZCkXOjc1LaZBiKxQnn1J8hDky/yqOAO75TrPKsCNl/6XUa
eKT7dK2iO0cxxzlSD64xQy5h9fBr7PS78VY/6Aj1HRbyKnMAXZh0rpJxwtbrAWiAEAYCA/ian2Tz
Uk+U3/AYOPhx6EfhaE22W6g1MxrPGczktoT4WYZ6Z4FgSzPHVU/hbclEWzjEDV7p3orGid46TWiZ
JL0tIXjlQup96/s+2U69JxdaHhPseapUw/inxPfwqTPTfrfDNR6yC7vLH712SCtKO/DaO4Ft3NCp
BvU3gUjbv1yZVp5QnR0QB5X01NSwqgIe5vKF/YzVg/AQuEgVowDnDyase29HNebkr1CV7Cg0Qvh+
+Hk3xKIn0EoO3s7GmtXGUu1quIaOkPsOAM7uEkcP/9i6jLxtW+QVQCneqmdfTIIEPpVh66CaRDod
VpJH1qP7Jduk2LT/JrGkpjOdAOV4g9w5OgstvL3TtNSmolDX3Qood45RtYBSY674apNRTGlkr65j
PrhfmqavH1bwRU20AoA75Lt2BbCGIUitV/NX92EABoqZ7QvmAswu3HZcOnsWBlL4G/vjy9XpeH5y
+xoM0u9aQXWLBpuWBDVsBv0e8jUL9LlWrfBFYh+I4VgkeSOoSWYN/1weBtyWd6xp63/mOwIpr1vy
X3eekzFbSObBTxKQGAsyh8UqWg7DXKYnFVNiBdB3nq3j2XjwhcqKDE6cRPcF9qK7HAGffmrSOcnj
TBM5xoNg9RQX5VLgZ8RB1Pq9nV2PLucxjpVnIzMV1MnIfP61DqoWs8UVzhVefxeTXCs4rJPGhfd/
fsSspvLhBCgxWJEbIRYfH/q+som+L2ztpEc1i7w5rajfNH4Ev/oJP6Pz3Cw8+CkKWmSNUNSkhxYj
skyzFaEpK0edZSYe/U41lU9oTz6iW9e/E+vpyehj4Suy6lPm7iXCEgjjuuT/5vV3KZ7QAg6FhRXO
bkvljUPRhoNpI1YTZeJNgIPYUGHsgdDOTHyK8U8gwdzudTMfsKOOpPeO3HftyL4mWkVIpSElYQlz
kxxeAoCMOyMZ1XKioknkxF0FOW5elmvjJBmvMJh54RYrHueYlyUcSdIzGqVX8Ez28CdHmf0fIbD5
a8/r6GQpKckxBImdekCQ7paOLtaKcg5W5B4arfLpJBzcY9n69CI/AViP6usLS02YMOUEF99U93C+
EFP04pgUfddSo0mKlLQx02SrxfRoEVYt1j+RvdLIsuKtk90U/w1vNBC+57x3KjOq2NwUti67aqUc
AoRx6HOnI1JENDReFYb6IYJtCNyRL83dqz4+3GGwyC1ep9oh8wXZ8zdyHmY8vyJ2fMRHqSgFunFu
TymTaievHnWoVuigj8eA1r3CSTh6+LIigr79s39U8hYEFQoZI88ZVFmydVzEqFjBj8WdtdR8Ed+6
t8x9zW6Q0ISL2bCvl7HbzsWrtRNCfyjdFnBN2rBilAo9VS/8/4X2sOLUqluy4RFSOu1Q5zPqN4mV
lVUMCZ5gSWAdYB0jyhuGXPVkGfBh8lZ3Yeih7qHG1ofUhNcraMFtLeShZe4q03cm4+kdMW7EyOO1
oSgDrDdCYsFHo7HvuczUNRjv1qI3e4pGwtO7DKJEC+KeRSkBE8k0fIC1QSfMJHvJg3T9VnIcIqQi
Y3sPsyKiSZ/s6VfqIz4bQ+qQg5m0toJ+lel72ngyHa8L9+OrUo3Dvw637Dk4e9AvXQ7eTB9kZMk0
FDk0+xyAeX8zJBVUFyVKdwIquKTGk1gsXFitTcnQjvp8hyIwMnYfBdKpsH9IGbIFd+bw+/zHdWc6
rmo6SUvfqFTMVH5FolqyK3LXK6pOzc9wSUuXrdaaqCnbxnF5QE+uknW3q+o24rWeKvHZDIpw+1bW
mPpnF1GE9wzfDE0asPvrRf4qokLWr+ZytiJvsHDXHxK9trel9pPhzwfmjo3VCjzXFDuZ73mb0fBm
A/AfdsxKi9uYb0lRLTot0cQI7xdB9kainc33DbMGkewnFnWmvdthIl8zNgickns8ftNfjgqppxxC
GJTDAKzvjrqO4bM5aGgOuLByodSuz82mBnVQqkEcKIIkm4NrOCJn5UJSxYDXiVLH9uEf4pqV0jL5
jzbdyE1ZU1QggU6Vje7Dv1osf1L4N6+/RmEs5d/vAwyG7XX4cSVtW5DHsT2sTQVL/RCGhKEoYm0C
ExwysTGLqykoX8LsvjoJuxMGYAZ0iu4828njnNe6p3oqyjzINYegMujtPLKULzeGKZEuvLPmYSix
ZK8tdevfObS6OIp4286Oi264R7POV5Gnadw24vs/m/ICUhI9Dyo3YseRgrON/XhPSS295QXPfHlL
lqCUCCjddPeb2h+dS54kb50PB4NOh9KopZ9IEngXOz7aV6nwliDAFMy76HCYJSw6OR5G6RZx9bf3
Oy4qXJlkMQ1QDBCZdSK9DU6mJ0ILY121DSDrZ7d2f+J9NM/F7DM51T+Foa/EJafQIO55nJSp6FIg
Pjm35K2LET+GZqvUfzODia7NucyJODTPBwlPHiYqTqJDu/gzMRWgorzuy9aQT9Sic5a+a0ysflt4
Owh8O7Fj41uOMI/TPrzqWv/r6IafnUY4DyP9pR4CQNk7E1VxkY6Hva1xi9E/hEtbtLqgZWwlnzgn
43axTo2y3iIucD1QpC0m9R8ISFQH/SPZVbC7XOVGR8KdYz+bgE4j6VTZPceB6r2083PATAMwGU2I
r0vqwl1/GRIUEA47o+V1EM7FwT+Cu90yJ2gWkpOgxEA87UOvgkMh3p5dlgQY2S71g7l/IxJAU5Ts
X/Sr+IMqmr8v2GqDqZNIyW+LPrKKUyVJg5WuxfDlPvyRcva1lgKfnYRC3gn7nps4vndRD43XpS43
5VYtfqs1oz392RFaywn3nVjsByeOq7YnofHOSgd+q5I0oZnYGqSMXGeTNxTlcRMlv60eucP33+DZ
hzsSpwOQ4AdzPmFTJebcXrh1WngFqEWRK1miB9YDeKbjS6KXeG2iWjK5ZUjCQp4dk7p/Vs+DNTXB
jdz+cBWyU38F7HNF9wxJJ/NhKLjPQfSUqFwsaMLH3TdB3nmj7IhJekopOjDSUO1YswqfSlXTC8V+
kouvqJd8NYRYvBKRBxvBxxFvgptnQA41Rzzqc/gQ2DM6XABEnOT0QvFXLjPk58j3sndFinTmAegt
FU1T2AFWbIVqLfvL6DwEBNkjMyqhQyikHW84CBA8mNGw7Gv6AlPmWz42zbj2mEz2oPchLTq7HOPG
5bHVV1/3B2IlCxshLYii4Pfo+IVbWJd66Hd6upntOmYoMN+l1iChoPGAf88siWffTYIDN44/L4ef
FbsrgeUUJLXqtBylxxAo89JJCxUM90D7gfxA1yTKPzP31hgW8QaP+Cd0Rmwo9xrNOIgq7lKSHCG4
Fm4rYFNQ4Q6qkbYPfB7WMFDUz7RhIQn30eMn5eXZLnB0dmomIgZwVnPDfDMo9xxCxpFfAKhXdTHB
SSbRQeF0kYMV4lu6jJsyU25yGKB2gZDGDnBYkp2lZcg12qY0BQNkkYiTjXU/mBpK43CmEr1NaLkB
HecuUjMWG6vrwjxprHxGyJjh7fOQk48sPENTU2ldC/HJfFATNuCYzP4IwNbNwu38K+Kf9cb+/sUS
/dhXQ/8Sg1PdDeGU1hWlUW0pn/VJI69UAjyCXt9bGnrgIfvXDqLlLBYMWwidmAr1P2lDNDPu43lj
kCKnTgaoxBz7+N7BpUs1dKQwGLRK3osY7unAg4WTABM/m9qS2h/atG5v3NAiVwvZ+9gkBNKUJVJ0
I3FOlkZnFrKVRdl/ZLR7T4c36ZCnYhrhEtTqXnCgyxY/Jmz9nwdEyZtUVSEs+w67f2LIxmKXSc2P
1IhrP94SJJQyc43MI0QL8O+Ee3E+YFq7M3WHQnSNk5ZNQgLZhBOc3RO7eDEd7B+GBKxB8nI+WbDZ
H5DMV5as6JPQQhwV2muPFJlLzyuInKN1wAeOGIWvWq0oQB0oL1KmY1KohNiXXO+9UXKTIhpIYnhO
G/HeLAOO4YvAH4IGBI+C3oCJDF9FPZJJycSGWBe5XgB+lDH19iu3LACn+rBdnenGN7fiDOe8Uagq
kGf6T30xyZvybb+YBU31ZGQiKVj/lePM8kUigxXrnCmshCGByH6ex+U0rNntgwLvPJGgzcv4udZD
B5sd2oLjZetD40g3DpbPI0vokagvyYnsYvBirzjZF3/U5hLp3D5+TGFiuFPqptwPcyzpnflUdGsF
YBW76MysHcY24+Fgu27iP8B4V7DI/u44lr3IfOA3MpzOTa8bIFtVfFPf1vgRT7+4dHV2wpMKxrHE
D6sGzmr1PXyr+VbPYbhfqqsiM2upPATrnASgOQPkoNG3ORpeCo2pDCVZzzWWq3gCKI5Dv5tfKWaD
C3qj0y6GhmGnlcO54kNJknSlhsgiMRfUPdxUqyfNxCKV0TAmCNWpjQsXR4tPcRHD0Wndrt2e+wHA
DRUZR53uLRZBvp5h/uzWyR77EVD5qmsQvcOwjxJKkKO+C1vT3+JrqjDZBAVMNuUnQPCvBDBOCRk0
PgR54Px6J+xfLug3AFEX+g32WECkL41/gb5I20Lgu+NBwgYQVfK4mK45HsHxAkz/IJXd98PX42yp
EVH8D9I2O8IPvFep2w3JXR3LU2XXHJadCbyoCOq3nRbZlV9RaCA30HHUYjl/XDN9cMaPjltXE9Lg
Y640Wa+TnooYpLII+bNr6M+cdasY1EU0t6wmE4RTQMn31C6EACOE2qfFAQpuEiZUhUvgjUBtxnUi
SVaXIUJXgAg/v0/VTaPfx17b0eaq+ZzKjxKH5mrT7OZDnSzEpprL0e2gdbJlpLxYzhsxkxdAJaVU
fCHmy//SEaG6bgP9slRFgBr9jg5B3CI1C1kkLwnijTwv7GuBcPxp2FSSmak28sk2DBsFl0835hUu
iMVMhi2KdV9zELmtJ28nY14E+VidLlsy9rMZrbQgGMocSfeDMAWRXrnqW0mz63/eI80COw2p98VE
pyWaBEOU3rP5c/TNMGBtDUNPi7CazFZvTEWOvAVIw4EpZ32JeS0DdRFzvcWJ/x6z54mdWx6xPBGL
Af/iCos0cQZO7DYsQrUt23Nc87NrjpRhW4P7u4tdwNnN/5hvwJhHeWnhk4gqsjc7ep4YKzKxpVHq
iXL9fNeCZ1P4/ya7GXsEuN5g9d/MZPDFNINSY52HLtKonGg0s8Sp0jxws3XFFNAqBYbqyssjqhLu
LrOnduUBa5kx10A1/zRtoH5dhMPh0JxrtW7G1jnsIfVJEOR7YcwkrFKG5Swn61GVY8zMSvlmC4DL
SJ7flad9JAWXuMa3MKiZzcec28LPjMSjHmw+9QUFKg7Jht3wkBe3wN63EmxRLEPoyDPWUZ02osnT
h153VvyKw7vTl4Xe3wtvi1MquYDBJaPaitB79noA6EEvq2oHb2DzrQRZIuPabuV4XunyUDNRCfe7
itmmz54jgjAt1VYyaWwV25p4Y2l1HXdhNXFSEt3CbIWHrGBnIS7zFvrapCoNq8UIJMdblWEc5xZN
ayVkUUJwJER+B0npdPXbm65vlp/prMJJ9mxxfHeekgHk90izWnT5GItueOIbXLfon7c5eTm5GVsX
LXFQCTuzClUqp6eK51dgo08EOR2iXLPOwE4LT1U9CURRLAWbDcqI63yMOke9VcahPGxxbqACZDsj
zNX+E5N6ZRZf76R/5qLm+2MW04BqYPjEBt07DsGJ5BCUMelYNlakydZb3yKktOi9dhuufCP3DSJI
4zNqoVunV4gPB3sSbFgkT1B/9Dg7F2OMkwYFzTarEe2MTPlcr8U1X1ZQUxDYEzjotNhDfKuGYbV8
SwOzlbsSktzZIhaO2ZVmSJvFSleqAkP2yKe+LylEBZF7fSgwHFB+zmIrXXPM7GGMpGXDXNkaWYiH
KHzoFq+aL1Z4HWE3zw/BYECP6wi1mmmdXDkgF/20dMgormC5bwQv4VTXLsII28Fr5YG7ja62Zq5F
ITmpx6HM6tCcaZlvHjnNUh9/iJycDalWtqU0+EbhF5Vg0z9NnrphyvZ8RTnzUavUgH2leaANUmQ5
3AUQ1VGZ4DpePDu0yJYT/Jdp9LZkcH/cwDEQB8CvP8Et6FMlSIB3V6KldMZHazud97+R69gcGkDB
vSDVnckqk+z8r9uwkVM8ti0hoP9eA5HXQNo+eoFOekcoDijZmJf/CjgH0yOkL8w7F6KY9jnnSUDd
9iomlIYeFEQYrI5ZFrpFDjNNDFm2KzGPeV04a2e+xi+P3qODhTkCmXVPNMlOJkWcNgBiL+1/twb8
+IS++Ygqx6eOhWTm+YFmoC1oc1E6h4qRT7TA9WUlcqgcPXR3wJ5D9J+VgpxZMx6bXsRdn3b96J4x
K/VYMmJAtKKAIoDwTjR/W38Dcqa4bL/I0ADi9hP26ddvVU6JL74mkY2iwKFbdlz8M96GZ3+5mX2K
JSJBgP6w/cwOQyC8TbPdZr6Jc9bdix5SwqOZ1HCArRSwq+BDrBWzb2m0C+gNbzptZy3a976c50g2
JEYR2x/rpJ6mIMNqhPd2aUPwQTEXJHBdTlnyLgERmLWrfU0IO4+jvzqN0AD20oZ6KO6x1zkRSZyL
TSXfGeLw59G78CmLiZjkaNaNcc8uzS8HLOUByAjyK2XywwoIGW3ZnXDB/7cAoOzkIBCxM0fnp2W/
4IDeLggen1lwsThvy0tyIPyB5XFi9GI9dehgHiJaAuUTYFIIbckz2Ch5CCmXRl5danN5/qZW3G2i
WIoh6rRkOBjU5ZgY8hMofjXeH0/3h/sou3/NPF52JlZNBMvWPeN/z2ABRGym5vGOtUqI8MfixWHM
MLdrvxqHgF0NSoc5hbmCDzpH2J32QeftS+spqc73C7VMrSi4ta24TuEQv5M4fbMbS6PMMnj4Q/x7
nQ4fjbKCswr+GuOyxLbqoSO5VPdYcRIBZVMKnk4e1k7vuIOrw3vzXOE5aCf3fDnVbZrXZchuVhZt
uW7XinC4uyE9ULZSX0m1CJwQIq+Kj2Se0REycn5eNK6ENsTsvM/Q794fg8VpNWZjB+vx9wB8UJfP
M9zgRIVjQJV416w+aLCnlqFerx0xN/aRYD4MOhIbeaIxh/7UJ424xqyXg8SPY2RorHjtBb0Dwgcr
B+pcg+lc7Uo9Y77LKrvcprKapfmVOPR2fgq+F6LSEn633MgJAi5sFTw+9BHAKMBH3rc1l0a8p55j
SdnoJsBfO5FSuOSIIEEkxOw4LmM8nUjAnTLI6ASld+Htz4hqmv7rCg9jTIrPYL/j3iVoxmO53Smf
Foye79A7ZssOTivbepkfQyh4GPpOUL7g994tcrBWmH/FEn/eXJtFeIa+OC9Nns1cywr6tESlnA5Q
jIGqdUANYAnVN5bnemiv2S+wdWAFQdHII9uoX6Uw5hzmWaGli8Sp8bDYnFR+Bxr7F88oem3iZwKu
7rwxA6Dqu8lc1xR7wsaFaDK4lgIFQAbp/uqI1sg9vMFeCmo6INXJagpNZ1peSuSPTWWIgFlpdsc8
1VsGAc7or5SfsbpPGJPdCffMYu0rGxjfIAX3KdfSeNYbI4y1Utje9lMW3y+WNJ4cUgZBBQP/DKV2
Bl13rsqE8hb+pw/IKitHu1NgsYgpVsebHPYj7Tlj/yyarhI/Kh2cBT6ZBcglcBso4bUwj/QU0Dp4
/I1ItlssAS8RJV647/lRdchfyDI3XxU/+0aqCi9921iyZtQm/zrBRIWc2+/2MsxHcJpLe28R752K
YVIf/48f5LJ/rMbJz3KlQYLF+8tvcRnDpwuVxn5Jy4vAzusTxIzXj9LAa/7HU5Lqx2gCt/XOR1Ms
sSFy1mTTdWh+KwIAFNUe4wCKa6N4/MCfMvsIpVDUz+AffgeCG1WvZgEfms7XKVUehl9Xzr6fFCkI
16wP7RuW/iDHhp99KXKXQZqAGH0+eSd1rlVvdm4SFEOHC2+Tb+rZORJ+GNR/88S609SeTI6cUvz4
JxjA4fspjHbBrT1j/tAVechI0r9o9sxm4kbfgacKMfCDBbJGjOoscj7bXNDZE3C+ZtvEyA6DJPxN
/soGVWQIZ+onMgtdvKORVSeBtvZ0a5Cgjn0zM7rGKyItXaSq/qJXOT0i6BRU5IqqGUyi1YJjabz/
6f1tei9DAT0EIcEkdCVJ22b8woAz7Ids44qTxnAP1nyo9iTMqitdMOK+/MKPNYnEPNVX2M3mhxe+
pkyeUV8+WwwrLeACJBuLh7Dqqy/p80ZLdmjNO87lCszdEzBwct1oBNeiPCuU6CfPQuAIHYUrg3r0
D01SaDy3iy4t2lcClgg8mLHmbcXKF6WHXp6aYl5YG8txvBpnIfhIgZQGOXQwOERCQyfEFOwOsXbs
wlUI9I5Aa7NjE43b9HldTseAc6QW9qv6iM5n5uuEAzIkSQxehix2uDfiXfuRMu1PReGoEDRgYe9b
huwASVOL5rt0Z5LtDd/nD3TbWQrn2UMatafx0wFPEB743MWaF0/xvdmeBHIR9GmxcZ1emf4IJI7J
1ClvkbXttFzXvaOYXw39WohepzfnuM4dkjB8fGDRMJN96rpgstaqfBkeXS1Tj+piojCsMw8Fkwbv
lgOsuQQvAnM7BOPpdrp9t26LwiLRZmavoAvauEeXe4dU+x/ypLSa70vqe79QB9Q7CYD3U7jLtqa5
7PaDd0jVKfxXVx/dsZzwLYi7mIQ7mMHSwjsHuVwDIkENZR+RjqXIIsnE8djvCdj1eSt3xJKxh/ic
5YJCb+a3osKM+oQ44wQnOSmSvTW0IT2+9G4u1TK1gkD9FAThp2kTnG1y8N1sB+Yp8AC01mxJ5MVx
ivcz+gpGHq8n9dMJ8FqWwp17LKwdAKRrMegj2nWIBG+t9nMXarkSH4MGPu1MxYDmEITdoCCm8vrd
rWLsahnsDPNQqtqFUeHgudxdGceQMHuf292D0ZSYaOwyo3W+SJPnyDTS8HVAjNwIElvn9hbo+IGF
XNF3ExV07orW2zjKRRxD398jAX4GCjdMzDdsQoDuPAy9GQaKKvbIk+CmVplW93OpYkRCK/NH2yf5
T56y1GB0XIF95eB67+BCM/JsbZIzWBCh0AFeiFiZbWMmE1++8JY0+nFfAXH1DEjOtG/o9HlbF0rM
z4t2pjLCKk+75Ts7AnVm2CPMyu/8M9lci8joS5JSihHLkrlk+QgXfINIzKGY/pw/3pRmV9yj1EBM
GBVIJPDL6rbb79m+D+yqw73TT9EI48ufpsHwLVKfj+GR1M2NfjoM4bHamJ5WRZo3SZGrtso/VA6J
cYWfSgYwXRqtAQ/0XScLTtadsyGPQ+TzK90YjZVmTiQ0L5gU12Ovls62VfqOiB6KtfNtCjW9sVFZ
6dxnM3pmJlR8Ei8wDR/R5zzsJPGcCoupi0RhD5XimUtjYtCr+ZOXadj1MHt2+iiHCppVmNaxCc+1
LAE2dQbUUAw1wxeRxT/K5ZZ/cg80WfD2lZb6N9YcPQSOHPh0djoWUnoZP3DBgJfHRzM1uwd6/2FN
YrOjzHOW+Wq+Z7n1oET+FX7f5VUNj6ovvbw7qqheryCzqqYpVshcarVPApKinM3RzBXnRSCtl1WU
zjm7BI7T177mNLGAamvRY1EamzBEE+ohq7YHB+rC5USIU3nlqDVgPmBeEFJDMQK5apBffe7RNISy
SVB8oxMsxFjHuzidDxkx4VCaMEI6nmX2mHugKnugcMP88f6oZKY4U3wGZJ5qRBG6x+ZGPn8XuKNG
R1e55H4tmBtFxze59VuSBC72ynDjZ6CjHx2p7F7WBzaJ1QZ4crmaB3/KFZ0T5nqEXd0aoRkEq97W
mZ0qn1LNdPgtT6I/R0CAMJeuD6DpYJhx/jT5eRz8Bd6J1H1eR5hhrfL5Pnt7HvKsz125lPKkAZnm
kCBOcC8znBVoxedU9jw/lkH4f0wGKnJU/B63OF3AY0tjFTuTRXCn+LmQUePcdYBqojJpxm0Ri6op
fBGL/0PYkeIblPo8dOX88ZqlnHTH9yYhMRsE4sSQLMqosVnJUtEO2GPnEVKszLp6oxwkP3IX4gWF
ZCbP6kSXgVn2VwGIx+JxKingCk67onwgI1elgqyN5MDUfCz8fxn3UMolZVXjgk0c/w+11XPOSX2q
9a6pfHj61F6UgjYIa0QOSu2UGZYUcuTOCeLFdqOClKp6y+QefTd+f4VNb0IXn//1oW9tFG8fF3hH
/bUhhHLDrU4XeHo2zNLl5TQbYm3fEyIn3vngkJjTCp8EyXFw6rgK/d99ok0/7E9vJw+KclgaUUnD
CiOnihoT5tBGgmPal25adAgn/pxLrFzRnbFWPi0FhDUtgiTLimY6anmbXgU8i/VtTPYoxOn0pvFh
oSJe0PsMdHbxEagTEY6KRU64+UFoNIZCWkbtznTzNjLCYRr2CZiM1DA6JbRr59jcOC56vth1IQYf
rROpo6PeSWefBhnu1qFAwJWKteLBPzYQ/X8/FDZStqVzFIkeNNFD0dWV8NCsYsK93PqiEhjS/jwS
GZLG3Sgp1PkoczInxACdkELmt0sbeFkMq5IIIxTGxeRdBD98YnTzqbtXNf5qLS6Wpkv/Jb1d1QCi
pFP7lQJpdcryhx2s+uVzbej0pegOfv3Ke4ZEh1RXUt97bC0AVQM1KUlU1DRSBz5PXbozeDg8vir3
/KVAZxiddbVHYJhrWzkd5F+u6cPl7BALNhFvqbE21vF4g4nbQPmYWIIkY40P8DRdZokyN1k1zq29
Oi4fcb4TBivzRlaC0E3M5LyVUFRBNZri2FvZSyyNprjVxGOHcH4fkJQcYsuWNrqaXkOa+J36ZtZw
7r6cW8QW0vmipbxHMptksZpqjYjcwHbFJG2kbDCxgB2/ein3MJ8h2x0avMv1qfQmJKs2f1YWVz7a
7pFmzKvXAjj0RW7gaols6g0YVa9MEqMzv7GdoVqKQJw56ac/47I7CxOqRCUMNi2tNr1Exgx6PncC
GLzrTOdigAK603chL69LWEBFHMcoK+3RHO37oUml3qHCOpt0omAtl+P70Q5idiyqMegRZZVhn26H
IOHj0lNDmEURB3ZlPewNePtXp2qy6eAeXvwlIlfbhNUkBBHnof2Fm/BBGA1L1k4w5FsokEjnt6H7
H9Ro9nvHzNScdcOdJleSeqcFjnUHILz0ZpyFpt12lUMQY6yYKbBDAalCLeHZ1bBp/nTOxwhe6YUu
FrEyWqMWFiYuIbbio2q5qw1FJJErk/oue2/Me4JlQvpqxLA66n6zIeFDhlXqsRd93JElBrcThGwH
q50m3ipcQCDUFeqIuiXvxW53N2fZYpIc/MlxPU/2vJUXJ9bYIUNS0G2BHq7KVKLP6wt1v7Da4NLF
4dyDLMJdZJof4Vtbfwb1QHmgQ9nQ+pwgLW6LErkR0pDLcGDL3EMbncUJs0c+i5Bef9eFIBuwm4Xc
/6FuKcOHzGQQkSDnpTMRgdp57RvaLNbq61jrk4DwyYoDygU7L8+yAqF7lsDn1lKrEjUPmzbQM16y
sLpUOGelRRTDvcL6G+i4xoFbtYtQvlnCLIj0E3ib9aYG0h52a1KRGBIgU3raS7fMDU9UCdiFYcg5
tVMyzep1e17cnHFj359bG5V/3hD65b0N+z6tqa7eMuRWr4QszPieA2EGT/nLR1agEG5AWMQ9vvB+
CrVhUQVbrDjnWWHzkI+h71B8sy1o+RLoXu0fzQ4cFFuhDzJQFhowj85jFqgffA25HsevUm4ZXI0p
vanjf3gkLi34blA25XEz+GzBVFYYCtUSucXVamIz9E+2Ik2AA5BcftgAfPfIBFLbSC3EoLpkGE3o
T0OiLiI2/bVEa9G6c4yhLCP1v0arxTSYUNhHSEoFBtH9hELKLNCMnow8He8MYa8QTNjSwkCHyfjF
cylGseXWc/bRHkRU3ffuijuW+vF9O8Mc+4SprMrJOtabxu8ey8dKzcIF/WtcbBwqlSi4eobU/8R3
7XZce4D1ES52uvPTlfDGUNUU24p0XI1ceDrm0f4zMl4H1YbFZL5SC+vPoFEJq36qiLoOu257Pc6A
ZUay3cb0rbx7PLgF1bVYEtaK6+uGyFLkJAaWyNpnknyOCj1m/T3B41ylh/LLJL8dQswbLmJhzil4
7o75m6IHSG+dhpGJ46Sr4Qk4xuHbgPP3XWsQcTDnzn2SO4vvYw433JmcAQQdmcPkxYPpdbQToUxF
+6B30Z3Js9zFUKl/v6EXXxQCcBa9U4AV1RTPEnnq9O+DjpTPY5yCraAzWxQyTBtdvisYDeVX+oZw
Yn5HEBe+8Q6t2eTtX14581ofK7YefhWoKo3XQBLyZKdNVJHxeBAueMtsBgFCHpyUoxo4DOTEunyT
Bg/AfMPiX8+CW09o6NzllnK5rizvi6R1k8sfJD2B42ADTSstSGDGGwh6ZKcFzCjBXfPbqtNsmLU0
ent4yzDTC85uzuaIUTAGl+QgZ39fwiuf9TYKitQh3ZbkVYH6ZZFbqxUNvCNwVYSOayqchkpqaHCY
Ryp2RpcIab40pBXMF/75PZowy3r8ygmwiLsFG8DjRdylD34kciGVEPYE6kaWn/8GsqAhMXN9OMk8
+9nKUtyy3UxQ82aJUC/Zu6RQDDvSPVWv3mr+IR8XzRjX7INLVykDUemx8Pay+iWWi+tDLwwrZ7on
f0AmeHtoX72SbHggBMhrdtRp8NrDD2/bFf7zSGrP/MGHJbwWLob2lszzmxbNaLhcMzA7cgzipIRm
Ao5LHDDQ+z6BfX5eNCEzNs7DodHv5SYf04V7lySqkKrSjfFAVTg+L9MCHo13qezgwz8MfPSVbKvp
qDR+dusn6z9KR6XR2+45/g/FDmhspUq0z+vuCNWD1lDd4uqrhftC4NV3MsB0w17L9FSdXhq3dgdd
Q3ETuLV63qWOrYjWh9601szUzFnbYlJY3qmy7QHzmdiYKs+megUCcvIhHOtMrblrek44We2F50/I
u/UNWbpyRMPiMGd1g0YooxvbeOerbMIFYc/WIH5tKTCzPmE+serDKdDiOVlnpIwv3slUVMUaXENY
WuKkHTYuv6rp5saf0ssJF7GOjGwU/FF15jTLdrfIVX5Tt/Il0npCSn0/w1kopzEA+5qBtHzB9cLu
PjFPZje9beqewiFR3pYj8iyjgdn3pzsakTuyEbvutsMgUr06WHqMDgQprlMvdW9n4FpB6DKvskg+
hCXHVXJ3/Tq6kMz4AMWkZPxfPwDZtxY6Ur7wGzqGsmMa3YTuy7c9yCr71Jd1V/6g7zWNZz2ielz9
VRnm7atLWvYTlPWUvw7Ur+ATv5tM0Q5ZeAvOXGchSOW06gq8d/DOr6JZHDoaZOIMRLnEJn03HWk9
cSfIT6xKr9xdICkOS+SXbDOsb2HCxitU6Y4fB06C78c/JsfxqR/RFukC/BvjN4b4DpSmmBrzBP/b
m82OcEZLCLpoZfCHGgPilp76kZtCDCOcOtMPPiGgt8PqUaBvD3zN0qC9sNJEz7xg8VrGvt7r+2v0
NkD0kwMu5bBX9HCL53SWfS3IGuiIT1Oy/Z0DH+XNMIEOL4S/eU3gMq27wXiqVKPTTK+wQWC6ET96
FfQHAOzyFL71mWm3ZGrbT0GRurvcREZBT7WnQjL6NGOdo09quMpiWH5ir83Uz4F6BWIDmEswCrBR
1kwK3l9BznS2Yrjrfh64Kx+gDyqrOX63261yv7ZZHrw7D2CIXb424LS02InUxdQPkjvwfo9+uZrt
oH7qNpIKeSXPvMPkrXxlYpMhnY3eWm/37VcOhSq5aETE7kuqVCkvYhUqZy+UQjvJN2FjRZsFe826
jWqGjkDjmcVNDYNloJTeHIsAhTkapPB/B932FbNxYemxVaPxS4BLKrP1eqyzkFGNuwnPHWLUCqnR
xVuEbhqF62MHv9hRKy92lHQbuofTWhbB92DmX5rIVPDq2YZ36cCQAZwCpykr33ivsmznoHZErS2h
G2K7Vk+qfRj37FEyq7GD2I1QihSI5HLIE75k9HjHDV2QlRcrXhZ/3/iHHE7va7mAqCUp1fahLNZ4
b0AXkQn1zhc9IItRcnEZXGVGzNXls/jImASDVbC3HHu6l10TP+rDRt9mE/0F/VDid78xFbV+dLxC
auMWWQf0Kc39hGmiQIq9mUKztsaeulImMSoM77MO1s2thOedqvkpoxRBKoQcAMLYdLSEWXKcmqLg
rvdNfkjaHr4kEkxq/SO9LASexroqaQ0mFI6CaUTOvNmhm6c3RI2SvIhjWEYpPRlS1OM1yQ/CM9EN
4uJs6CmopRLv7MX5GaRMAHkLGgs44Aet6yVgXeUkpQhFucD5YrUlF5LubdCcIcjGFD9VpMk5eqnF
Dmby4Zik011nfR3ihbrq1ugJiXUFeZGL0BGLqTdOWGsnykISydbciAzPUEkVIch+rHMCB/V19zfk
iIYRqa16VfeEwkovVbgB5YwkSRgC4pNIN1M0Wt7Fmu7hDapmPlzHPXsSC/ikPz39Z9KcfanSKms9
1kQpwz/7aiQKKKWOb7A95iRj6x7nS/vJNPm231XqIhB5sjexVTuJ3lWE0jWGMVHd1prIODF6ltMp
de7xE1qBgEzpFq5Dv5V1q15/erjUJLXyfORcDpBicXKyQoNuA8zL3rJpYLBlhAmJYZaKAKkI8LEb
cquAhNqd0ZSWGsqiOk0LqE8mJl8XRt9xH049a7do7XsHeGyHWspGy7qhRE4Kw3YjaaLJJfhWRCua
o9CCmTxE69T6mF4Q9qutptyif2wZDrJPxrtjt4HBj5hK+2FreHZcdkB0w679PxXN8/lRYL6U/khi
Cil7EWZtWyB4HXS8oQ8GaKf5MFV6m2DssVAMs2s9UcWOjEX5iVRcwGMa5CA0YmaIJFEO+8jUSTU9
udn3hbkkZHnzeLFF/Xi93Zqf78CeOWsDBG98GUFKPYNsHnaLSHWl5+9WmvT9HdeXY41h0/j8edzG
OjFE9BuioyBAogRiH0GQl7KALBP2iK+nXRvCWbgE3z9qwHUBbarpxBJq9n711NOlHOuk30U9SF2x
zg4oYKrtyYqMJ7ndXiPRv8aHyF0z97Xpdwgh8cDkIsfi/tcgb7/kxzZ5OmA5xWVx6LYgeTdOUqpk
X25PbTI8zBT4BXaDMt/dKNrsWDuZIpYFJgHY1VBqPXo0z7gsi+ArIhw9IkD+5sfmg3VdZGA7ykve
cQuSO22q8f/QEjcF8GABZuzEJDO3idcaoQ4dFOGdQ8gugPQbhibQ740mu0YQeyVmOVtvGXGgi2RP
dANA9IgBGiP54JKcY79xkm2itru+9geb9R+Bj3rk2ldF2Cl0DHP1hSC1A+8woRGKsTkvbDrA1X6z
1gteGvKjbH+/bGhDM3PYL0wWXkABqR0qhPCFX1FK0EjVSlNi6z3JtfM77Qa+CKZIm2RXPynVQ0Bs
yOrqL9R4Av5tZHVe9gK6mTy57/PmZxTKuQaxcIDJkyFtNL1zayLSggmMu8JjorqTrz5OoKKcMtfL
+viHa8vICM1hgvoiIJy5n6mTB+ZyLeHW4UGTqjTMY8MGfhOGiz9oVLBYjFdgRPXXP+GJWhC7Vwag
omjAFje+qVg59iJmZvpLfkW2WA7K0+FY56ap2bzEfP2eTx619QJoNqrvLzOPoKSsHsJF7s5NYcqL
8SkiiPkQ334qSsIFGaR/978gDiVIxJ/oQhR/5eX6cQyr73gLoTwGyXApwHVtf7WZazSjAwX97qSl
wshJZU491UWETE7h0G5ytEIKRxi7nhu07ily3r5sPFbD1cblV+ohNPxTOyT/Z3KVpp7y42VMbzgr
mcFW4emO9ryAeNZfo+m3vq5fuJRwvEVoMB7ATRjOi237C8ShdW67YBePPObz4IKLv9TS/zvQyuVe
MHTut+lKom+B6O8ECsK06cu0Ld18SZo+hZIn21RcY0de1zS9HUKDeAalfrsOHdgTZ4i2U+kzwf2E
VZmNafo2sgFW5ELhMUFszC+TJyn/MSQcxe7O0yQkOWkQokp+SOEcq33evL8y0svi39h0fsqr0LFB
dMyX/qlMkUuiPOBv2x843A+7qHbkTQTRNr9CLeY0fXDlfBFeKJ/GTi2do8NE14HOyMa+i6W6PWYR
OXTqT7oMjmsPTvb1it3pf7twoTnAIMzzkW3gXJRzL2q7IPTxgY+t6SJkrciRmozalUfQWMgka2QU
ytuexp9AyC+rODXNVqatXXEsPxhDtLBgHcxgadAEfGvLG5WbZmmaNL6k/rT4pkSMs8+afpEWixpV
HBYi/5HswyQZwbktDrcQ/SCEullK9MRsaxdXJ0UM/m2b1nfQXtIyN6J02j74RLclaMJ/juukRdfD
WHI0OVwxhH8l2MBuk1IuYK/Kt76jXgKueW2Ho3OjK6BqV45q/aam0v8nKDEtD8jItKMvOhxmQ6ZU
gvpri0MmBaeQRnx94ej3bg3OkMTmEfZgXflHjSQ1G6dw5lSX6wRijCpJLr4zT0fQokv9wQ1k7CmM
Rlj1/LI6/iz8Mhsvz284t9yWbQn8UZCEARvjEc8go2D0Wo5M7/wz0FSLkp+YWW0XBqzfH4X3kop3
1dX01i0yV7bod5AOKveT+FzTxmiAxRaNwniU98+t7ZvdbIvPVKmHqr0atLwqvMhVknli8c5CZg0W
CRYw19PUstm8bJLj4c+tncGnE9TVYmty4DD4lC3ijSSetI0GyOwwqrilQRCJ3KiUb5vxu7ia4wFM
QgUkesbmzCLZzNUiUWwqOWrDOyX6J0vxhdLIbpaKJNAzx527fPQFK9b0/6S+17p16RHCTFNJUh5Q
asppXe29jYAEJA0NcL2+MCx2pWs17l/g4jQsSoOVMqEdwibpK2aEebNx/LN1LVgop1OfaR+gob8E
bRCueISZb5HAc3zPfHq0fOOMZOWzqvZcy2WCZ1x/aFYD1l1Rskd5V52YNjfBo7gTqRBw7Wd7dJdC
n4WT22wm16utObtr2W5gDgUAzHMJqNOZdYBQeXkcKSw5uvqPtcGurBHsX9NWJ2x6Pd9wfmGLb5Yd
+w3Aiep+EruJUdVZNEjNeibDL29T9vch9vtQSSrgD8rV4h6dbs1lLpXJNe/MseNyOIeVfCcA2oby
ZaR1JQKGaQJyHnHGilCLcSF6Ngzv3OagwTq5Obz/hwsSu6vhr44QwuY51GEwwg7f1Y9lSmyOd3Vh
r7z6ijlmrR7BfgxOV6pR8vYbV8sbdV2bQXU4J/vsJUOAYHCiebrhiWaLF32JGLv4IKijhTQf670V
L3xt7hNDUAPxE6lPZTiMfAALUpRFcgtk8WV+v6lswQb2xlJRvbISqwmkkdPrlR2hlev0gMZztRqm
6kLhNa6jnj+SaFJqTRoaxb0xGmInJYi/dzGbzNBHO7pjCZojC4BpN9qZLHwuglGnTCPobO6dA/3s
eHk0fiKlNorQbukOAhe+s+Wpnx/dS30/ihCD3sizett0XsKMoHbXCyxRnjEOLhxtjRC0fzE6TVzF
ivYQnl2nvpsOpGPJZtTQwZSaSObO6aYZnViZNNr/IRoeOuPrSF7a6fhubw49VP2ubiTFXGf0pm9M
JWPrVQpyyF9GChBsRpq+SEq6QU6q6wsSDwUzgfSWagyQQGiB9UOsrSZFkHYUKl8cPRRpCSR5bws0
b3xqOIWvepLjJjsATkzbB5l9Yr3WBZA36f6KVmJ5FgDKCenXSsqCpwrvC7qURG/kLzcNjeHpN1kX
JtpV8N2bj8cjrwMldSitqFjLNZFZ+EfV8FmL6jeb/hMkZFH+kZWFe/xJ7iqf3R6V/9G7VW8dtUiM
8XqvsOSM4/p5l8p03Ybkb1le4NlcATY/Wr+/3yoodtHHzbWNfoxkwrKwD6TvULMH10stuc3VcK/u
cH06IsGqQNdiEbfzj1OAeBKB7MLOXe1Tc+6evfyEvXsXQrcDx3UVm9oV+hoXPor55cFgnnG0BNnS
q88meltueNd6gg6KSa71qw7LTyjAUDMMRTw35rryz7w9nQSayMF3Gy0VYfEGD2HhbNwjPg6nprWY
mx9aPqQ843QQvRZB1l+sRi+scIgPdSRhS/vxkV1AVZHGkspCR6cLqO95wI4SSQ0BwPafLhEB7QW0
CpHtG/42gOw41PPOEDa50K3Lh93ltqOvSiq18ziAORqFTAqSYKclO8FfYxo1inpQxjnsErR1U5SY
A4pahdWj02e2gSKbpYvZG+EIFejtUDkSWC5kblaHpTk08hBn4CblhLYWdW+QHZhVxnacIfqWQW4M
6L3mULEMkMOcKkCyzuSQLcvYs9EHJ+OvOLFhaA0OdEzhKChURtHbPavB14erI+lrbGyfQ6hWd0Zr
+Bb1pCMgJQSNdeAdbJ6WikosRy5ypMEOT0KYwSADNnVBLbv9GNHoqzrh0mFuk1o8oD58alWLFO9N
wIOH4rv4vTXj+jym7TGhU326nlmUIfue2AGD5qynkupShUYD5Ld7ENo9tRvF24QvcGj/xczDOv8L
05kb3/eS949TU+xMdns0rlcSPb33vCzSVH6T/gXQ8fxAJoffrlyVMaBTbjceg8WhaCZbbgeNsbYq
pBh8PnAtr96Wp7tbf0MlchTjzO3NYvw8PqErHOoO2ks8G4vJArIDjdkmNsasTZ+z4Zc887ju7iJ6
1qrmew24q+rlT05YLGfX53kOIiOklJyaWIzXQneYW55i+lxixb4kuBzSleuOBE5meBTXsfIWssAA
s5SaIKr52c72XeU0hQxlTXavhnuQEwVrNV7XnAI7Tshff/nyvMAb2Mcnd438J6+vVXDfKsuTrAFw
QqCbqvIn6lBi57Db5/ayNbqukKAHlZTiLBsuB1pzD5aAcShmw9CHOC5DPFSwC4pVx6OTURL6QZYV
jH8OaV4CRMnIYvjKJaQJ2Ts8IygCUU2SG6M2J5TjM1r92WGvR9F41k7g5pX7dsD94vUc3HJQnj4C
KokQI6RIrGQ/U+mdkm2VMKe3ESoqdtnG19ffx4jhEoSfvAlU5GJQ51/yHouTb1rTMZ+R4cUuvPx3
mSCQigER76SbY3lD2Zwq/ccgNJzGJbocYqdQDYO1ElT/2zHswDfeo1u7ymelD10Bq7iHoXrmPriZ
HasHNL58cy1jFbfOqUrd+mf25sgfMJ5Gvtyh3nqkQEFoNw5qNi2iqI2svnCmIO3BlnBlTyX8UW4y
DRZ0yXIDMU6d1UJedekIWYd7c2LZ4eAytWkNUDdKMnsLFQjaR71RJxyDjPCYRsn0HF8lXLNizXfq
bFcZ49ALjRem5Axy5nWIkeOYXn6jlzgW+ggHvUsViaoLwSihjNYZ+NiWr8FwSzpfcHmPxZEvq8zZ
L7OwcOZZry2ozIqqTzRASr3dP0eghDIdkEVueAAhpCKhAyGU9TEA07SBHM6N4+gIgdfP8Vpok4A8
BwtclSHw1v8o9WrPBjIiixfij59C71IEq3j6TUAP9yLOYefD7qB9J7mA4bsm0pG17Ny9NttPzq3E
NPXSV45KSs6rjuV0P2myD00p4iDgqEhTpBGtoU/Klw3z4KHF4K45YqHJvrVBOeChRYkmUD4THGZc
gK4bPV6Hce8MHzX1+KNsw6R641mv9ilU41nLqnJSuysYo9ogoCo0Tq1T3pS0QgHjul0doW/DV3Pn
cewCDvVj+IuZ/pmLKvW0Vxxf799rBmXeorUoTxZMbz2Wotse0T7JLx4yUVryw5zAZ3R7dUndrn/M
Z0Sk301A2dqBVRPXOwnlizyVlZogd4LIC0FDiAWSgyt+HaPkD9ZNGMQKYYYbxiIx6qRZJ+KG14T8
sk5AQDmivE70V7uMfKeuZb/ggPL0alUc2XEfTfnhJ+z4KRgDHz0rr53aZmvQhzWU0yTaa+aVr2ZR
Hj9P6uCwF2Za+qpu4vqWi8wAkMHRxZyMWhyRJNi7WcwnZrsK0rmPqyJ/5MD+2CSzXO2+YREdjBei
EUhaTKw6mGRJXmak6cwhInt8nmtKVwzfVeSPiWyp0eSKtjtGKBpjrAXD9z8ijG6f0/xRSaU+l53g
+FcJiFoHgl9DSmpSbZpMn3igyS720lW9A6VPOXI2qWdoJ2E2cCzItdYr1KRvNVa41Kj6dJJn+lr0
jygB4Rhwp1M2US5GScL9Z4iZkWz7GOl8hxk2tUyAB6Q3EGy56Bdm/14rG6EWFQBCmjyoN2sdhcf7
qiZIJn8LzXftTUuQvSQ9SeP+NINjvOldNfNO4nxNRz1KIrAC7L9Y78zIjUf/HsnHd0kZwE8tpD2w
VKazNYweEVkwNV7h/R3YJwZUMovjDjPnIHPww67BUzHU+9z0yljY4MXZfsaVux2eTbjPpktGg3ua
KhObM5HWGBpMKSTi4mJC7zbl3u6xMT2k6cKMFjRpHlVXa5rTi4ib1N1BjM5aGehXMoEg/D901Ehr
JygPm+nZwiLG08GABijbDhA6VUj5eXIv1D+TFGz9RyQVufBd0Yeok7iRd+ifgGiL9bIIf1Z4g9f2
rl7luJxVOOLZv7UkMhA1YVI6Obt1JfluB1MrSyTYdGGOY8QNCtuGvuHl9Y1FEmAU6P/xW07imvtB
+9HiQ4pjjFtNaHjWEUFPQsKoFxVj/pG6nLECADXuJv9hUcrRy7f2b5EhDVW/VNqueFQuAfCIB0WV
jdCmSsN4i+8wtM+RIWj53x9TV3SBmmuAUAUjyvFSEXrKBB1QHwWo8jwTTb1PyWYvl9nXSkwUZNkX
YAS6615ilML9lNfH6pcOXNk2Xyk/T7yLpLO89uDlG1AFrFMOTk+9W7mILjprxXQdFRs2i5c0cA2M
AlFPufvEPqlIvKxK34uhl+FI7ZIMLgRLEjHw+eE9gyHOhq7ZaCi9OGolC+SnXhBO6UfY/VJ4FMsJ
GbX/7/ZAj6YpBEUoNgEWUuLXS9ZYu4Af5TZSem/NClA/SklMggvN0NZzJaXPu00/RNwIVQ8LL8Ke
uNpqc3eaCcFBJ2t0h7I2egiidffEIHWFeFajgsitsC04WUzRFwY7GdOOxBP3ZDuiHVI7sUKKMqdh
n18wVCUAezQtmcQLSs4wvVavWH2Kkx7dwdCFlM1Vj8yZgpbW9YuVHH6ErQnqmZKW5o1PrJi7L37j
BWclOPaV+5HrSYUvwzvDAoK307tLmniDibMKNc0TGYjPosPf3fpmAWGSVQKl+biRDuu43X1VQVT+
s/qUMjSu5YU4rkhiTw9mW+j+mOdEsaRgc+va0NNbHB7jLPhHE+E9/+QsB1zZxPu5oxJas2Wk+CWi
S67H+flhfTWpc5hxan27RlZiTLxABEhIz3HgLGU8xr6X1/KH8Vz6cRqInxEaQ00MtlL5OunS6eA9
sNHGhjwrcsNEciJuerWyqPv8xlEkdvGa80I1TrUOC7RvL3xnlhQCatufdt1SwR19xnxl1rM6xjqm
gpItMmztOI7CvMLvgmLiH06ehjRIPJLH09MlZ1Pp9tqcRV8EYIphJPjv1nZZiXlEUZSgs0jUhMb6
pP8GqzM+zXBA+AUM4TxIoxSboZfz2XaEmjvJ1GAdeqgYlc1K+hcfVRBivEMyOfUyVEG5MS2R4onZ
SP17uEVz1KB0yv4Zhvd1fYvBmPXRDSGLDe19qppW8NXKqK354cMQdZtb8eKLGoEZZg0lrmTYncjB
rCgnAt44ueKDQHTUZKqvRqAC1A+nlL+KM4jLO+RMrQcgBzTbcWYGdG5x/yIUXxiFWON0e7qS84iR
Lr78TQ10sUPWCUbstiu7vrtNc8ZfQaMOTyc6yo0bh+KJb3UTGaJBMah5xaB2b9ONPS5ArVbw2xf9
Tykz9wg61HaXPY4CtRcsD5Tac2i10dRFAppkp0TSG8kXVxVEDNFqqdCtVhLEzKyOQyuTuK+Xe/N1
nvXKxsuFDmF9RnBixQ+rvS8pckieVOW+0nYMeHkUrDt29lXVBX6KibagfUsm8bAt0LddPJVrw1CQ
mCk/PRJF/IYKe+7phe8FdObky01QejYOsFxOzqTjz17W59Op927Qaxn2uXNGPJfnW2BHCS8bRjcN
BhjlRP0ZhV2MKtH3QN6K5vsfkSg9znJiORq7vC8ymKO1FCime6Qs13mpH2x88uJZLbDEERhn9tbg
kbMFjEP/MM2vtfSIFDmkRUhMGt67t1R0TogRwszW4f1SNGHgzo3CeiU3GCBug9SEYxjvqOg4IPfl
+77AyJ6i8McxZzVoi0ixCVm6uaoKtTHBkINXakQWGojx4VpVKYH8dHd4LW3ZIuLncR9eeAnqw6HL
UMj9jmQItAe87XEpUFoEioHnH9LT10+m4rBUz0X2gVzYS/oIYfEgSL0iLJuRA/V28cioyEuX+51l
Q+WbeRFlRCgLzX9/TVsFNAdxlByhaI4LATuF69Gx4bVsKoLG8m+z1M5nEYPcrZqfVjSA7tYp48D3
wJTNPsENassKLbZwyzqzu+1JdbRfFChb8yux1OLnBrxSKUsGgkFyaZwOBk5U2ner0B1OYKCDIRGf
1YYyI3o5vrxnm1LWkNZ4YAXzYSNrB41tnsIOFLZKk8v48rvTp5BU2gZ4O7GG85zztzyPzIX7Wsko
JNMWbgcbWMcWfGT4r1DOnKvTKq6JGB4waa8YngV+GkdLRFE9b3kF24WJV4+YR8UJVaWxdlZk0+Df
SzBsFEsuKYFkN2+dR5JS9SaKJyEWnbMaJD+8cMPc4ADE/DmBxEN3Tapx/1fTjI3lDz3Yd3ComzyT
R3uMVnDY7hFK6wGaRFua9Htl0lAoUzBuc+Sf4kcmT3KsCyE78I6AJemQESd6l+qDcmLG4Vb3IB0I
24ZZccyRszHywZFNB2eQCo9QxYDkaCSGoG2fmdI+uccTXs1etvigVcGfXxn3EFigTTBmWEEyXGyC
nKhvewZbw5ZXsXKv9+ofLk5Q9ekO6EIiRDolKQKTrUCY3lMvMzWHV4471GnTPevbbjE/kraY2G9l
yBGs7j5xgGp7aEZBwpcbzyxPM2LBTzVrW97RBYQddgFnLTws6hXlw8y2LlwO5fcovD8roHWU6z+r
SEttdFnze/A8xb4g9CIoJGjRpvLLCseCyVx71wQZz0VzEQdv+1d1/3+ENBstqIRHWdTkNdmwk9Ld
dI1i+5uPdRi3fVzrbsyPemUWJ3OjFJc3CcpTRf5KACn/tlBgfN1oWdrLu5ArtsFiRYubkbErZnBQ
/vQqzBNvjHQT0vIEOgScyVwqfXbTjYArzu0XvmSSLIujbl80mW5x7R+pGBENZY64pWjWxkGknOxX
Y81wQAT4soQf1a5T+Ddj5hY5emAEy/9Ke4h8p6sjlhkEEGZkIePTli4zB592fstI2WR97eUMyUww
k8OXbs1irufT6nxtH7P8I6Yb9iDXt42eEFOh9Dl6443rYRwsyqwXP2kyTKQfSIXaBwwqVLkZr+HF
O4mYWCmu2DwdZd/o7m1JDuEN9DKfRD497CNLXWp+j3N78QnvtjmCr0uUAwoeBgGzdyKjDSuSvy1y
USod+LyA/JINHvNQp8C1/8MmhKgx7qez1rGmGzHgxj2koVeFBzaP2I9VJICzluegewNuXL8LTrYJ
Af5ueH5Jc3F02opi9dnMN+HN8xSjXIOQq/2av3RA4dV4fq59mYaVU0NdM5nl45+LEivjBK/qb48/
eCBDyunZSah52HF0KyIzfUiN5O0Sa6zkmU0ob8hDp1POVdD4R2s2ltXSNM0uEAupGHLoFrTKiXmm
wfR2PXvnxojGFWoOZA2MEv0XIJu2hzjcChAK2oQA8HKmQr4CyTn1KwS+lc4pyNIpl/AGtBS0wDeC
xWJXjvoVoFrCWSsuaQaJLowO5IUrofhksOynRDezI0PqYcCNyTkCMtiCUVFU4FtIuP7l2UbYGs/Q
7Vdcred7gBNgUfWlar6wK2RRbylv23AGrxZqEyCOF6wusbYcoOSRJG1/In9en9BNzKN97Vh6ysOm
mzhjEUjIqkNYf4X6KsT+4RVwGN9fy4ydEU+8fqpyv0sOpS7asvqGEOPgKS8nluSYizngTEKxSXD+
dU6zftIedSjTEIV/88QD1BvfAmelIBOCzrIr31WTnnAujR6HmxPMl1S7jYAvw9mhP5+yWD4Boulu
6phmRSNp9XlPXiveIvz2L9AYhLxgc/YVM/jlN+MxXxQnsuMENrOw7VlK/0SFSpi2Q3giIrL7LuUR
Cd0O7mxKm/Z1qeN83QmFRO23VFgwSdEifYXmSNkKlfMOoENv6TSIAdbyt393funLF23fCZD/iVPp
vo8NgmmlmUvDhwNgDfS2wSpo79+CTHdaspBSONRqFUCZPZwh6YJtTf0KtpqiHK0eHjFzBPx7C9Jd
/sz17jQ7qzpTP3Kq+ZDOmA7qmajj0yWXmfKF/hj8S/sPRT+36obJQLWt0k858xbHRQ9s4yfCOHx3
Qh6S16hqjHcD7Ef6I3K/FIr5fUi6st0MK9fRD6Jzf8cXSmcU4Zn2g8uVwBKENcFCtlOxHHtAhGrg
JquHCKzysxvbvsAUcoar7ZzgrttZpO9i0f4vcfDOoeHPhZ2oRA29qtgRnE2mCwIWM76wfywh5RXi
le/URD6m44E9B+Wjyz2xELKhjfxW1nhmRYylKOcssMWRxhgcYnKb4LX0XfWsgaCAaDkiSDfZ9Dc8
4RvekoOduj2cTDw27S8ziEUZT3gQ3QyDbhoKEFKsaX89LXiTIhKZIaYabFVvSJ20gxEq1BtILJvL
X2VWnZIpUfsXtOzqolmr/PxGwH1F7qJ62c1c5+PWlFqbS+QbXF+ANmNkTBQpaqwtDFQ2Z89pWlVP
r0v/Vdc3NfXRND4gUnMci/CJUXQ30mOc3HrprfPFv1XN4Af9/ZA8/9oOpsLPFKLyeWE81O661DZa
+CCQZIyhcC9ps1EXOkKjTCNg50BhuU1cxhHGVMv1UBidNyu+jof/nR61Q1DyR/V2/dfh0NTa4+rx
g0PsTnbEJzlPX2TfQ++rfWLFFnjewoTJPBvsxO/D8X9pwkjJdhF6d44Wxkfahi43G26vzHuHULbc
+vyQ4KAQyFNfIPTuaiTsKXUGJVJXlVwna3PE00ySUAIyFaVLu93XmR3eLdO+eAfum9xUXVh34qam
adfiNJO3biJpFEX3CoqhhC+AzcUg4AJZstzgL53GDGd4Wj7itqU8rKO6kyT1Ib6/ZBRaj6zK4w1m
cydiJQGPs/ir/cxpdPr03g4xZeXss2/gxisg6+qeyE0+6JJqU3HqYfP0jVwWVlsBe66g9c5AUFFA
0zAhNBuL7gZZ2/YsAd+KnpqIroxWHOE7rgeiyP2IwcoHGIwaTsjDShJrq7xZxEyk54SJKaAMVSal
Qyp0mN3lrysQ1hX4lJg7fKrNOuWu2dMKNWiGYkz1JtTUAslw1Mm4XgIPDJ//KxlRD/No6I850kIn
DhkQ5bzS+zo+30Ko57YEnKgc2imOPJ6GiEuog0ghFhZMLG5E8t7I/qsGgoN/tGnDmYEDjWQIYDTk
gppdgSxAIqfEo9mRx9yTNsQ6x5hUcDYiGMe4mefQNy+PL47PQdmsRkXirNaHbdhMeOBwFPyK2sqD
D+fhVzB/N0t0laYcBkXCb/VDAwnWW5IJR/SrZdmvsbAegMzQls/5aGeu1SWWnYKBLD5sD/T3W07l
GiiNiaupBapHUqgWJHJeBX8wAuykLgN28aecY+5RZ993fJeYAMzsLwShkxDNFskyrxO/cqzmxd87
PdBmpdhWcVRVPtoU7rZaFihfWi4peR6oJs1kuGgU/iYTGWxuItmR4KSZwef9p0Eu7VLckIGOTLQx
BzKElmQPcvsXgQWpyz/+2skTAg6E8gGtkoN+g2m9LHBvPyf52q8e27YbhKYJhcJGsswlrpheFrGk
BGryP3pZKJEC80rRtc+paorMj6C9CdCzm/6dfniv9BKlxCuMBgVNCPYqfuIqGp7DCWqZ3P0gp/ll
+yghvAO5FpKjE6nGZHbVkaQrl1kYSJXoWxlcmG3W56ZHqRCD9jOENoQLxwvgVpHJLHJpXM210bU2
99n+Jwh4A+hUJ1pRILeS+KqY/AHAheT+6Hyu7CJ7js+jMqvja6E0N0BZf3+F7LHVqU+NfXKBYdpa
RTyYi+T1ez/gIgfHR81vha1eoBM5DUYSAfM8FdVGZOsmEjRd4NhET3x74IqS1xAOYMe6ir8uKJ19
EWs2KwsjyhfBkEP4yInyN4D4GFL5CIK6MriBVE6cf8MyYbJ5lY6wJC8PNGkO+6eLs4u7dzLYVCDy
J+h68OO0ciF3SKF1vtuwgr6dFpUmC1FjQoctmwxLbItMsyeNTApXP0nqvWTOu69s6b6bzD69fI9W
z53d8+AH/JswfqdhR1zjlriuyEfAAsynkWkrgv6dZ/MAltGAoiQId+7lweUvlHMcMsgIfu9WS0Ku
M3mQ1AMQA2XgLSgG+f3Emj8K/vu6gWhW6Pzl86hGij2iV1axqIp0c0kenoEaF6hcH/+W0oQ1rNe7
b8HLQeWCxAjVZexJDLHmb6HNOlLSSV091RyRW+4WsM39jdwvczDVzmarMYRddcRaVaWeHBBBTrUj
5YMObkxgwOUWZmPw/UugkKJgqopHKv25NxLArl27XWLn0D2B1YQvTLy/eP8xqK4Mn1HhZ3rD6kr4
OZO4251OL0T7612oK3rQmKpEd7dKA6vr0awjB2bCeR8mGYhgTwJAECW99eR/u2ch/RGcJNlwXd14
ZLSmNSQGGJpYWZCwXTGMJHb9PoEIxc4b4NnfGU/cUsUM4igLkGQjJlIPzMU7Zu0L+k7Tr4fwo7k0
e+c5F9EcjWMSIZgzGPjF+gOaUuvOHU/3iPxOpxtqOsi3y/N2Fc1XRvZ8Gzvzy4+6Jcndfacql+Hp
t1LL5wchFQ9xKy00OpoKbgxi6VOPTPiFyzMG3e3nLFBwbqD4hmHronTHqj9wk3FLNxTU8KYEOJGU
wCXkd76Yh1og64JPYK4vOhF1lTII1szlXCeuVtzRbyi6P0gGk+UDRqwZEK6Q15sWgSD3kCiKLgKe
6ouF+Lx39Vya8AQJEpFRHyvUlc4brsfWqnZuVq0MF+V4KtDmtlnMTaLMfDbP1bGsMsfLWOwJ4be4
+PH8vdHSjPZ3f/2AVvVPQ6cBtC38pn1zMtBlzOQhzx45rTDjmcInAaIwaNTZvAxCCzklJV2VWXpw
+SOjj4j/AqOwKfVETKo3lNRWdj8UKuTTW/I1zL12cW4iDs9CTQTZQCx0z65qi/qBBCYArT5Jwx3C
anMZdMX3LFkseb1b42v9zLl9IVl40V32EbmIwcYtjrO5vXPiQnRFbITePRB/JFbfvvDWruz5GGvV
Lg14cfHssLdSUMFz4CwI1OfpoBM6y8Auief+dk5/jzLe1chMVisnb5wyqcdf3YH+0NWSkx28unMB
meOtHgI5pAq8NpdHdxjkkIAh+6TVGf4l8AihfJriiDvuAe62HKN8b/xMYyXDrCrV3MOXURBUQSvm
0Znknvw6mp86WbUTIQa+a+025DcjmL6JaE6AD09sVBaCvB/SHpKfOlFzOg+Lte6OHGOyKL+m5MO3
ZbGbPUAbewgFLlj4caISNb9PPtPSUOq85nEB/VvbIA5eVGzUoiehHyj4UGzJQM9g/5HzPEu4EDjS
bThQ5jLsk1gXK3dXl8R3ibfEN6dgQfqw+nmD0/A5IBDlMdBRHBknero75TmqKakDQkBLzzxQoiKC
WG0xqT9kHZHx4FJ+EXN3yE42dL6cgK8BOi0OJnv/kzZ8x4bH/L4oRsfkMr7B5B/4MjXE6d6eugpu
yurIuur8OoJ2F/zuszbX/Aunm07u+Jfp8D9LeM5CVbe2ERZBva9e6mjqP5uVg/yIiohpFf9ix7Kq
EN/qeKNrs4c3ixBErcM+R05KrtGM+VMIPNys7A9lurLoiXXOXwHAZ9FqyrYS4EBzGpaOFj1Z4Qn1
iPrBGRsqgsWk7oVuwaXMao9NiF4iqcrPK1M0Zxbm52qQK9NRFMjsyY8DdEHXU0Z1JcJqFFgt5bB4
ZzWj/SYUiJBQTPm5pkhQ935agtCnxDev93d8Qmg5FSW+EYri6xjM20xt6KxwmbpD7RaFfpcIE/pz
7gbQpui0i5cSaVrNNTZgSC/fJhZqa3JfEaEnFwiX3N3gvX4DIPzuKa4twH8nimfLjMCqfSlaP7WR
+DW+x8+LQIEAbpo+q+G82qt7ii3MxC0AOMo7INSyNibuB1UnJqcycjp1euWJMnLVgxjlv4Saee8H
Aa6HTRBvxAoBHYl6Mo70vIkeCEWpTfpnWXwm694sP2d88BNn6cCcybS46rh/c4jOx0Zh09thUib7
/j38GtnaHGgtlwXQ4zfAUmkab9O1anQSd9ZT3jIzaNupZbkazu0YK07zLfBq5FeVok5fN8K50U02
MU+9TEW0sV3oQOq8MSpo6Qyq8UqQ0rvRLG8TJuKQ+bjUaCx+T3DfNPASBdxyKSwB6c4EdJFpirjO
cY9iungAXp8APGOI5WX/QMqggdMjBR1dMXsSIQKDYaeGHyZIzha4hScvpJ23n5nAETaGbwjbPgu8
aaE2Z7RvlQSLLo9YMHfCQFRXR8DqQK4OSBPsHB5whnC6dEBkhBEmXWI6hxP0F8ouS1ht+L9NFv82
DuGEVOJWT8HFycDNe8jPdI1iwelv+gln8hdRq6OSlOA/z/5q7EwsU4EDTmb0wqwafgZzRTVjyTl+
LTkagDm5OQ/EMxOR9dsKcuQqZXsXWMt3l/K8vjMi7KCbKcWt3cppKFD7+U6nP1PNLZS7NFRGwfXf
7Y6HiXthfds7qbCvGwr5//br6AnYbFZJu262lSxya/slHeJJAExfj9nWxpX15Tm38O1rF/KCSjkS
UPF0zEfcBtZq3QERPsPg/OUgneRmDGIgjEZTDPCeEnQ+760mNQq6+OX3RLmt8e6IV58PBq7AnZiJ
BAQuhUrdlzftjbQRnHsVWYY0lnpMq/e+g9QP03VU75kFHltZTfzQpri3k1AOHyoyuBuyAi8EHDT4
FCfIPvghN84M25pQm1f5+kscM6IuFRScefFy8AQu7GcpnI6Kxw1/YrMZuSfQAz9AFwN09sAaeVI7
P7PpS0tro4aPkbuECNU0k5nVdlNxcQDoTHSfyfnYXQC8gXiwoBACqTPSmexChq8BQ+EinsG1GdLB
Fdf0ycvsA6vOjDcRkrFAf1O+6IOeTNUqWgAGM+vt8r4OqwcwtdkYeB3rcnmecnBVLh8ZUayH2BVt
U8K4izvQsb0Xk5yd6JpZECEQZLyG4DQ/51FQc91bkqDsDEqMHpKBuAz3MTM3CY7f2XyUHrZFv4bu
K0JviSvBnCFNtQy7vduub8qGNQDQUqo4aWWXFgVRiSs5KFmTHCuEOkub2/FqP/atAWf3gh7mJ1zc
1ZLfu/I6sSy/JD/2tugUlgMj2wNavPSlqOFDdlMbDKQc2EXexGGiuSZaoeV/1A5YH7nczCshiuxD
exVmA/pcrEMd5keBzdqhcbBzBtKeL6aKcLxFZVhIHvLg5cbD6hYliUxEuDnrTgDfxxR3LDt3EyN+
nwAXgNkzGqJwwDlKkGAIrYxjOOtCZl+81XdFq5l9EVlanmi0zq6U/nbFCM2y6t2opU7tcxgHEC9W
7wLRfzIW0K+PyWB7M3ienGkU1IhShepPGeGD/eb+8a3XsfmePfo7yfKcsyHpGnALb5paa8uxlioj
OfvU7eLiTIqQPxrajadPoPKQH+ybQbPVX8ngctztjCdpX1W/dX/Nb4/ULF4tlK/ZLNfM7EBA47V1
5FgdDcn63Lys+QUV3cmd63DUk32ieiahzXT57uNKRmMAVY7gXIIjmJc+bh7g2aH1aayTuD+Wyt+b
lAbBWZuVPSxnrbG+n9FInrUvOWukR7O8hhlRkYV2uRucESzHY/Zlkf88S4StHnGI7gx1w6hDckIV
+FYwWxtgow42bqTojshzyNUjTCN370ddBnv2SmjHXFTKUc31kFsQxTXESyndV2gSMQReB/CuyhjN
ym7sJ1/14DXeUUHgjtktweqXlTsSKBs1kKFiJFyNoJf7Eoq4wVBrjJ8gs9/eGlKjdy0rBCP3DGIU
C0ukVDxI5/58W1lmhAnskug2isWy+2OGeHd8pCWvJW0Z1IndziVBo2P3E4/9Gg0svpf5W/DMwFWF
d3Eh3QRQ8ADvx6u0aWZ/j/l2UyrxhRq3ehRkU2nkg/6P/KRYGqfnlZuoi5VT/1CmlTg/oVZ41bMf
TGRCuPFmBSPlH/g4lO/FdeFZcyQaHFd9fOZ7ZwN5RROHAff0U7dVTlEUAcUKCjfJCRkll4R/Kz3B
LONEpBYRkcvbRtd5tfElkau++sfzowp+EjXgE7iTOACm3Cu0q6jG1qFkg1XJ0rF4RmldiaQlwjxO
3fVwsOWB0fz7TBKsZGVRLImgi6aing5Xjgr/rCbbTJbpgkEL+/0gwf4YGBjNXpMg75UCHBRr0TJR
mLZ70aTi6rlSPIMAECaS68iXwIHnihXmK5J0mdw0aKOLyoppEH3t/IcOr1Fd7V83lQXjInYr5nGc
CusjK9m7rCsdGY0XWwg6oeQxT74lD3UNHMPpKxBxRUQGXg6VfERkqsQYXvrLM6dtKCL+r09n1xiK
H+z5x5Kcy7SD9hEqrpPlezOs+vGw6R0VvNUI98WWA/cxLOclitdyRxPWo05kpqwKNcFpZbj6eedu
ytVXvJSh/sJQtlcZHSjYglLIB3zID2n+pP9gwA11HkSEUqemqByDTJudfENVqmwmWVAH81ztg9jg
SA3wzx2PfvkrLhuaXu/7eBWl6YGBj2W9VDMR/iUBRFT5AIS78gbpR3LZfFlqfJhkv3ApAShYrFI6
glO244+dTDxxa4xd66vCK+TOJIWdFboC9FQXNo7p3w7K7ptqGDGfiuDKlp6z1GuU9kPbp1uk+BTy
Snhf/Y989g7+EiRDg5t7SMdK2DhF1xtI642yqmDk7iqzp7p45Fgk6K7rlyHItZs2AnxjcAZbPbMC
kMGgwpzAFxphn5U5paYi21fE4m3vdWuH4oZXZui+KkUBvxbCGEgnf76jc7NLpIdZFEwxiKktg/dF
U7+qOrZslyN2O9ORxG6rVL94nSABbE2yUF2A4khcTr8DIbYt5eV+vNtDupQrOxAzXf2UXqg5gt0f
hEmK8bFJa97GScjMhnTT8g6Ch/kmMRw/8pngl31Xcof//4hlpyZ0vxSH9FxIM/7becMNbmJqnZkP
h2GMZIF5Elfcx7HJBqrhASBWptJg2tSYAE3SUT2WhZD5P7PXp5gSMb+i1wr45qTODn1kGxT1KfVK
ZRgwrhT3DjkTRUmXPWKPRFBBaRmyHpiw3aLZtWAgY+EYhxdI/oRG58pKQM6KPVzpfaDb4gtdw8Ct
GydSYfTuTa2/Wvhbc7ENT5KDUJDkayBM4zoE8PhCfI9AjSG4rbFI/wmnohZsOrn4P8Vxcenj9S9I
HILaMKSxKGZy73ZZDz1CpNZHNJkyBzbP4BSYUF/1tRRI0zGhBAfPz4M40EoAToZVUG6J2J/x6RIN
99bc1B8Xuk1q0G4c5Q0cu09V2CLh9ZWY5bOeVC+L2/3VSvQ0+u491CztYUzMdmXEELEhwGSx7dxZ
k760XPZhSL2eRbs0M0wgbOjca/j2/j3tiaeoD/bsPlI5pbR3+uTvLFq9FEWe5KZ8NSUIbAvjknaw
OZzyIZlBNcNJ5vRNI2HIIOxZAs+lJLoBzgheVJXZMkGr5zxzqgFq6AQ5NlECsOCOjiMMLtemacWw
Mc7WCKgDQNHTmuCtMCXgI/LsidXwXPFdjUt+CaNOqTQhx1sHRXescWBPF2S66+RZ7OmzCizr+XPA
LyR/na4akKzxC2vcBbflaUQrytStzOFLpdhXYTospi9Lh09UqfMmEEpe4qvax4c44K5hQEvsa9iC
H28+Msyr6z5laJJ32R5tbBUYhn+O4/O+tdVywnhBmv897UAC3s+X5wISw+94j5Le5bvql7+g+IGC
lztM24x3SnK2pgGng1Mw0Gj3+a+fTAW7r2xmfjhGw4NNJQ4F2KGW0BF1X3nlfKksC/hQCgeIDYE/
ZqJeUiIbYyO910BP6NoRG3cMIHaElMDt2O2HW1TGmwBh241QVTD5KiktzJjOzPZLp6lt3oDILKXu
kaH4lsIQeHN1WUb+gDrthj23fV3EdQC8t4NgZ6L2SI0IQ2zS66R/0dRPLSnAbRfGheUqkyE7cAvT
1JQyq5JklEzo+up7A5VQ5kgEAHzBxNsJmaWA7R0oRXVwVOWmGVrxS/PI/4yG5hPXbBxQWeODzG04
6ZuiHSYF5W29R8lXtEVXVsA/fF8tw0zDGgnhu9ZiRyzzaABdCHw470WuJHHbPn+gDrdMW2/zJUm5
3YJwGwAYIA05npCY2KEnxVXLKWxCaff59tCl6NyrndgswvCHH9A+beBH56Mb45Vbb0TdtKndz3J6
i+uL/kX6SmDMCxlMY2W/ukUtM6+7sDmmWDiC6kYeIdLaWEzMB1c9IZVPV2+eVq7ZDagyt1DzXfkx
V0M/tjNKbVS7WwL4FdZ4WywTTED7hXNDBzjMGOcZmzdjLACOtiqi8qxuDcy6sh8o0XRqv8a8QyHw
cGC5dqDd2WXt9N4jdhZkgXLlAIEU1mpvbuH8+KIOJhWb1DxOxq+19kO/Npe5WOQHdC1Y5d2bRMWB
OW1OnUAAqVFtql14Y+KlvNJnFzPFI8htv8OZlS7yCyq2zuVIUJA4OPlyr82I9fdSCeN83/Kja4HD
aSwts6WMOS4kjA1a4Qx03GbBxdN6YQmUA5Ib6neAxQ0c5Vovc/qBSjLo+5KUUOKitNHdt68sLxfi
QURTXvOoEhmz5kGI1DqWT17RN6frPmCaIPiG7iSMIKQvjKjAH0MeVQojw+m/7D7JQsnw/wMGytmK
uILsTePkgvZEI1ZodhwFbprZZVY7oZbXDyc0WsqRS9FPNYJ+Er0iP3cRRfMckJFa0dAN0jgOvLbg
+JwBVGdPJ/F/umGEkXTBNzwZ7chCx8OlCr3HLFxgvry0NhmYfNG8krYDWL7Ogh0cVzrLEuQEebo/
PsNz8SP3BBYCIYj+ZzYn1o55pcREQqiC8oj4Wks/aTchvCdDCavQlfYXaZYy5EKsX+Z26FtLYNOV
s3ipdR0MzM5qPb76dBheB8keWD8EInV/C92nLib5n5jvNhKIdfBb7E8w5oY8m47Nlt6MtUrOVzuY
vrUlquNjNENW3HSZYkPB/KZNnDmOZkh7j9dorbq/MBYLRY+mnRE9WFI0FfN7ikaNL4w7AtvAL7l9
wMA3bsrx4TM6QcOOO3dSc45jtbofL8Hu4qMpwMFpWchOF7YgliKeGBKUQR518RUt2fESk3YNmkA2
4kvNWzD2Xhf+Z2tjVuXuPRn4tb6paKeglfAxIuGAcbpyj5CrUVDwnvmEeIuu/JdfXDJWcM05bQhz
S+GbXIf/AY2ir99vV47EsSGRGt28LDmfKGbtOyhdBFEwj4x+/tPNaACptOj0Vc219kXhdrHgw40u
UfCpn3zyMFdla6HB+DNfpS+3YhwYS3mp1ls1z5fptcWTVPCHDZDOgL1/N86e+1jlP2m+fWMKvQRA
kn0yevhoUGrCtXMnPqMSP0J4YepMnhyfybR9zERbIWOzC3JCN1imZGkDqysg3mEMgLkc1QNBTZUk
uadYMLX436EmvHDdV61nWK5h37tBBfM9xuU85EWcPP8BDOdLnftoWfUwdlHy3nHVzyDluT3YOFaI
sANtBCi3A4/LulQlbzbm/oJWEZww0442/KE/wqaNXkJyhhsfo1Ro2I5zGfJjvvlnnVa7pW25e75K
UKHetSfarTMuhz/JylM4au60x1AFjh723Bi0Eu3TP4xKIiCGwXea8GGRhdsoj+dkT34RMG9LVnxr
GUCitLjl0mR2eAiOw7rq2EUqRzbNanNxKf0YTyYDVhtROtSgMwMD3iUKmHPIAqKeN7Fl97x8+/jf
k72Xv8dTmXE59GVUhB/MzHlAz41ScHiG+S9EytnkMRHmHMZP4kOJND9bmi4crhUYr2VquLzJIox5
LqiOIKmMFWpIydtklEevlOiA46F9ZLmHFWqxYKbDsvkiLB4xDGzUYn7nCFVKaDPTwHqSevJ9Fs+a
dXhgVp4esXMRRVMwwcj68RTA8eeY1sFzDHLihexNUtPMpd8zmZExOn7Kbl4srBhEe00r/OUPOosP
CqhL0XNLkcC/NyrGtux1Bb9JnjF+brE7D2NafZCSs8xB9sf3Dk5DxUztgguQ5YtPrZajl4YrEeQl
+xU9CuX9Q7sw+Dnj7QKZqUvzHghsdTIWVNpKCuWcGT2w/1yxNBevGbn06Jj5+v9zUP5KKZgMtZ0K
i9IdmSj394cGfM+pqtugrT/SIltnpahr8sYXOfcVdOAeBqJe7qH9RecIYqcF6SU60m5sevgUmuyL
C2lQAaig3KzAIA05RGVOlljHdy4P2qWyLaDqA4hHppad7I+9C2QRkKMD7qPKa98KPIOorCefeKbB
0qd262vr6CYypx+S8MQQP5H03HV3p4hDUx6joTP/FirBFxUthlyfWnV27EZsgmTbwhMz5e2Sk3i8
kuU3jnd5GckZBsaQX0aKACc6P58asqgvGPJ8hx1lQuJ0mhn2zTYN9V3OOm79J1GHVogXJIKnbmjt
BpSFG88vMKRuDHxH210h2opWKncumlX+HrxbwDHWYEHfTQZoLlSsDgVDOI5yRPFD2kmb3vcULfOF
vNN0TQ1W3PVa5R99gZXs/AN5iYWXWnErXO/63Wb3EZzDeGWcM8R+Bqftobfg9wNgLVDxmDqku04K
Xqcet7XnbLeor5tfKvFbuSAVWOcMwMjDXdHOg2basQfuJZ1fwt0R/HlL7e0rbswLRy/1T098j5RB
Vf98qFPqSA+BofiazOV6HGyEwR8OfYk4CWrnagMUTPKxJ+FBEeoYIwoBZ4BuAVMiOThVu/fCk1If
30KYhjjEBlmrpT71UKuL03nx6Dj4tkKnZr6tNfjcje8nZHNxRFvbr18bagepsAlrwzlK2KEfRtnc
Q3bDM8brd7B4cWCQ6oFJedU6+CANYXIqaBWGeb0+EDiBfGUodTLmriu6TGpDPVgfDq6mAC6i1dUn
nWKU9AtY0puzCqbdUcpRJQd2Xc9ql2bTimcZVBWW0hytVVflcrodmCwcIw1CqCr0+i9b9h0WTa8A
o00GjozlH7Vm6hNQN2DshRNHx9h0nlzplXSIUmDJ8Nlmf0ZgbTM0t73YV6iE3739OXTjQmDxWHM9
XdsXHDiuhuQo47QJqqp/F6J/O6Tmi4OLNjU8n9fa/C2f01+Q5A7us7GYCKaYxFTRlDx7ilyPxHJo
QpzUMJTPYZyp6mAZXA+I5A5vdrYpKlVFPi+Pca2DCEjn+X7MoGRbkyuKQ9KVpJpnt8n0cUZk3UUt
n13zzM7p5LGLtLAJH8h3TEnp3jlE8lhEI7phPMQqrJC0vlKWhG33OmzVxVDUn93p51Bf5ii+LI6M
/qQwUnLOAfPB0h16I7Mt0lcnLDggCm80keIzJ+BhpJK8GNh84wntJ4nrsnALDhp1KR9YedR1OCSS
CH9xGRzrfrybYYI194mN4x5CXXAsqXXnN958aJu4SlSco+7pNOYR+iF0Fc6Mog2ORHGpg72RbFYo
U6WqhBg5ijyiWKep1O2+9wWn88F3830jWrG4D2lNuqAFJPcuIyvh5kzTA1aWoawNGKm0HtWn9FP+
zD6XjH6gJGn0zMnpPaAx3BDNPFgwaoHckG3aYVyNl26XffjpPy1QXAb95Owkry4eqMVZfV7QcCnb
+6xLrVXB9AM1aFuE/ep2+k+YzBbgFVk/HTCx4t0vPt2ildOcMMhvXv3fvusoHzCksa0Gl6FXYhoB
JdyrCtvgWxqPgcyaePau1eoHfRSZTflBoWwxqlaUSpqLAOGghZQynn4wXo3r9qV8rwioPvQJ/Msr
chwiEqQgKgoCCwgV4S/+hJBW/NcjrBd6oaauxB3Np94mdUWmaRRB63qWBuRbr0DtOm2XhhJee03M
BYId20/ZHfvcC5LS8y53QrTacPrBisWsnAKWHeM/CVLFyeQ6jqlszFy7dkuKI8/+FIOsRDnr/M/n
ETc7YHTW4rfAcoJBa0ui+kiRbSbRggES5c9t8stGSYCFKV2GOJQYxQIV1OoIo7t3iaGljfxUjxQ5
AIyJdw8z2dloTnBft4bBfobyWOvJ6I/cIO/XWmAudHD6aaFqFBU9NR3wWmZLuYsaD6gR4JmeLZuD
fA7XyAeM4Cj2eyy+hhJA/k0QWAMGj58XQ9AdFSi01fT6uPWG9gIrlbFTQVlPUk4uN+DsxzNwE6MJ
lN0jzYuZexE0sY8hemRCgCAEfmd2xKYv2YhNcD1TyYkcgxBk2qloK3i5zKn3Qyd4X8NdGZgM5T6b
3mh6lqL0c+rvwtEubRa4Qo6KECyrtXQ4//7JtKmQc10Xa/HnFdUqtMblHdnI1AlXgOxlWoMI/Elz
bN8Jv9wLiCAu5SzQ33CVbgJlrm6NIoXItlPzIZ1MuSrSz+Dfs7I44UoaDMCY0kS6csj7oizJEhQV
o40JsdzLrPjo9DGY5czdakruQslU6vKAqM6dD3NOeaQhKgaE2RBQLvH59ekPhIDC5woDalo4CUHP
tM7qv6/1IVwTpMUXywkaVdYLc2fhmG0dQYoFhKrUICwJ8+ey7ZJNoGyV/I4f1G9wkeI+dXYplpWP
QJxQmXO+LDTKJU28hBIT3nGW7p13lxOaRekL6F/OJJrIIT1UZBJ3NOsnKAlXF/RzVCn211CT+O3Z
w6DPLjAZ5zcDhVdiQ3SGWKEbc//hrSiF07cbAd76Y8QcbM6KHIY9YCC2rZRQsBq+MD7qlUIMFyY3
KbhQDiQ/6ofv4UJQk1UUOda4SYQ88aVaDnjz69r/t4aezY8g+rk+Jr5QSsOuZrryLuV5nTC00YMX
RR1kzkFdKfLKJiUGRuhd/XpVx+39C/UiDRRpByooVWNOlY55PntxElhEnxHjPpOsvY6u2c8V4sbY
37b+yUMzlO+3FGVawToEWF3mIeAhut8TrQYoAE+ILCp/WNXzyFnXi881TDqVg5vLD0a/tfvL9/ql
jwYBKvna530+iy/fvkf38Y+2vU4GDfFh8WOYBHH3rQrEDTT04hUo6AWmsDHms96QATRau1GEjPZy
9wYGvkRxL51nPuvuGiuZZBS0/iH5/VdZbBro/XboYqblQi8R5PLhP92wsYyp0egtmtQ5XwCfhjE/
vUo50Mex6Mg/g9pd+H+89d8RzvMAJKZJ3MQnAvlNvSucIt1MAB+fUR05Z2u/1Bs8tHjgGBQULuNK
BmpdmruQPk8Qifm1Xf2tjpwxaCxPxyRcBVi13aRwaI2LUkUhdSBOjiPPPNpJjsUYdw4mkfku97Qg
xg02tExv/rAIs6irnzMMiqPwj7aDrB1rd/sWkzRt3Gca8rJb0xzqmm/8FguZGIbeQ6avjplz9WYI
d0Cp6bgHoOVhxcv8pQDVyQxWZzJ1Yx0vMX6ojzZDnAkGs0512YE2zjv/Ozfpljxx26mHkaDBNRmq
bgNLEaDNluCOze7Jcm7kDt1ESPBoRCaacCmX87EKCgOzUfbIY97ztGbFmwSMIn9vY7QfThouLg9C
ZcecK2EJbA6B/eTDWezRHZKABYoek0rRdpArikJeIwemm22J9NjRSdk/g27Z+kIwLnz4fE6MCkUk
vtdyIQZy+XuAnN0Z/5xdPUZiWfipfhelFdfwyYWrpUob/CLicyE29ocCfmgKssVxgl2ODtSIXZJG
R+EWVwVOrQ47AgYsKVnWh8NZvt71w1chCjKYP2V2TccTCCJywisxN17AFAhLwHqiljoleRkAsagu
XIIvBLx+AqKGcHsfnT3hMJy5Xb6+r2kbDjVOlUl+RsUW8S68ZGyNqIsd/f7USXUxAs7+TMUdtUEd
9jJE1xFTRJc1Ug+rUm3QjKU0ppIaSKiL0WdwpmCRWGEuahC9pYf7E1Dmx+A9wSAy6eKzv8Fhtrw0
oKyoUMt4CtNVnC2QEMzfpUPZEVaspsIYhxVYXUd8XLEdx7QzL9HaDBTSxFwFcgh7gJR+NhbBYqXv
b6UF2JxDFK2NSyug/vUXZIyhLxp6z5p2QKo8blskpa5LOgt9yAyW2liSTfzmJqjmGKx12/wJm8eU
ugZOfw7Hd+Ww+DrUxP4r0XiqChkLllpKxp8ktXRfGR0mL1cekncpFK+QCV/lE08hJCH1E9xdwf6y
tQWGvOJVtUlTK7pNbR9pcYnYHoaHCqst1w2hi5U/wQo4WRtRYZ7qxfvOxR7me314ZmLHzAPujQmt
ksGMkp0wKC6EXaPVdJMuTCTPyD9mTm8CjuQIhLb26iC3nD2dvu9GlD9pWdWEC5eVQ0piHCoiMz2X
t/3kBaC39qZEPrQcZ2in/aF+KasOMQfOCZeMzvAYXpvBrfJtveS5ak/k7Tf/bqsg4QTcx6c0nq0U
ZDbEf3KTo52+tmJp1TvmcdO725fyRl7cT6q4ar/f7+DH3gIfbNMQfzSO4SnAAUCINmZepqAxUHhJ
xQd/QE/bnYZtnbMyC/OnJn53ytXRFyvFpFEJRhydCc0GBJmCK74re5fBhoJPLrCM4uPnxcB6xqyV
iLUz02oGLNRMmmL9zSndjPk9oGk3fR+2G0fg36C299LV4M3fLaV4Q+eJieP2XkkXwoAFpGWhYtKx
QQ12RykX+lKU68MsZNHn/TYx1H9QfQRFy4vVpGVc0TIEqgPKEoo2BemP6C2nb6YzaIquuPQ5mEKa
uDNC/PrcsUkWWQ6ovo2EmKM/BpzN+tjRNOh/moUFHxQSWx4zry4fr+GqaMo675OeTKQ23dZKPpNy
Y7GPYDg/rR3ucAfk4wtvS5JYwtFIRYfI8dQhYb+zv0dNOxHEIzBsN1Zy+do9qURdWrE0MjAmrKlJ
Es3Jsb+TNL9wHXcGF/GGfQXIjP0RRfNeRTkHpxNPCHVJhXpRh2gCq2KuPP/UU6W9z3z4K+dBBl8P
MG5Aw8qSOyzZN4lDPiRp6nEVAAUuPudalPGJ2n7NVLB20p2x1P08uFczgsOLT190LsmhkJ7AiNVG
hFUx+5ZUxi5yfiaYWxeZuNGEPEJIN23vYH1yAGGrk9mRhaZ0ec3qE07xG9U7UvbRc97bLUJVWqSr
zV5GSb2GpZR17orN0QFpTOpFRrlQmBN+AcYpIRkZGEJMyqIxGUH36pa2eLKE8JcdhU2SfI4Ao1/3
K3ueRfMSdMXmO3Z6Tq/Va4/ENnyVy7yhguuTr0KVc/MY5MdaxUyejNO6nqcSHe/W+S+yV5jAbyRv
JSAXAUB2fpRJfEjMFjgk0YPLnZ+sG3FylSx/GyiteovK8XVCsaVA8ASQcixe9ctZaglDaL2/vJ8d
RRXCW+DVHWOxPXcgjFFunnNm3rpADadCLgXYk2yYMwX+4aoImNqPhZQITVAYLlL0LiOELqkF3w5e
2GTQLvqWQsiOjHsDvRdbv7bFndAxdLl6lLJkKNXdoBXk9jhFccPPYfMsKzLmhzFmW/kz8pGrjfaj
HwW1IbO70lOszlzAHcnpQnlCrWNLZdDM1mcq9cCdcLKc/HLFUWcIMn4rgQaLaRpXRZ3x/KZO0Oh+
sqNCaXRrc0ex75mt+z1d5DyWSYCy9HF6IZdN290amgEAMU+oZSjCwg0QCut4Bvq/Dw6+IUImCazx
SJxy8xPnYBHQNxzHs0QFg20q0bWKRiKOCYnuVky1VsqF0wL0WecGE8J6LdCTa7qUHPtUNfRpuamq
acOYD3JfV0l6NYG2gBCALSF1sNJgBrwzzMXgsFrz0yfm56yPB/YiyuT2ry2d4Y3zD8X2TfTV+4D9
dWnrBJ1bYOBWepxvDFhtc0w9w1ZN5Md3c7PLcHnXJ9uhgrCxjwqXhmce1IbXBUIDi5xKlzIVuZol
fFToLmufntDwZNkdmKsCfCtOm30luBZFZ4wysMAgYUEB+40RY3QARBRrd8r8NXtJcOUmNjFGDp1T
BN2x2wdUj4/dy7Faw18AWpKJJj3Fz9e4Ki0TRu4k4VIsGBtvHIfcqi7PzoCqQ9+8U16u1Tp/Gq20
kfemBfcmXdgRn/HtP8zL49rd4/CxFZ3mooadriEea0CRDJgJ9lMvkjepKeoLQBmzi8lfSOsmYHQu
pWnQm+9Spq1kc7CzHOVIeqe7nWL2KJP763R450CQosm6kstDO0LPJ/3GIkENl37rNYCK9fp1c9AN
9R18AFPjTlzmytsnQ5tjW64KwrPZIiMgfzopwvVxvYV9QgtjIC/JBD2bqqsnNNt4qe2TbzG99kq+
FE1OAGlw0OkmO28eenmrB3sYsej8YDHxP9DkHIbSJVdL87D6jKO4PpuQwsNGakn+kf1t6PuN6z9Z
USbyDAanI1boOnBHD83hzYZQHNv0UIV6ZAf0oJakCv8croWdLSBQXAQGFR6MD6awQyKsqHpHkgYo
6XqVdSEJevMw7EyQE6CFNmeKm1kjZD72X1CedpY7d+cLAN7w/Sd0i+bZR1Rv7JJYReBBxqoP6fGB
0MjP9wT5eumdPwBvhgRRB+NubtGO2QdXwLtpCzz8SFfOtu/r8Gm6iC65jO2ZhgASH/GEh5opfokV
MM5TzhPtsqNjl/coTu7VEKERBIDFB7G4ZRM2YMczdMLVzD9tIRrEtWTYbuob/tEMexrX8g/99IPy
q86KjGxwyyUdAGFiCzfiqSEGD9c53IzwmvDnDN1DrcIYw4huSErZGMtLPIBd1ETy5mQoaOqanICb
ax25TjsMWsP2/g5FVds6U1qQmsylZJGEEr3ct4MRcgbIib1QJ8PFkVVao5ygdE+ebuFpz+tuYlH/
vXjMvEl/PGIf492Eb7XG+fPNedWD76vdT56F3AjoJQABVZQwmUU+CKT4oIoFeTCWOAf+YZcUFJqG
U6JDRZ0F1ol3omAnfXODTlfQYbYzLB2sgh5gs5ETfJKN5ckq1R0llwaJXU8ecVANgqPWSuunlLiK
2sRYe6KTWRoq5zXdTqTkL8cnRDZdYiKQ1b6jUx+dYCoPzTvCkYmZEuOyE4DGkMXZGFkr2maapCOR
AQVVlGab2+zbHXp8eD61DB7Bk3JKSLZZJOAHzIfT6YpJRJIwbtu7VA+ddXAILQ2Lb2u1keyRfASi
uxd6ajV0wty/bp0oct+dSHUTMHB4s+6vtMarg9y8+V3kwqDj53cw6skf+LgpwwHJfAk73ISAy6/c
4vGhHgWIKu3e4zznbXLcm6NcH98siCU6Q84yHUCKnCdo7Gm5KzmBDFnMZQSyED417OLE+vxnsf7e
nCSgsbHvZM5FnOaxkFNgl4pqcq1h+ZJdKXCcZ1sQVRDeYMAzTgv+4+wLS/yTJnkIyJKiEfqCRXzt
Q+0vPjSgEIzy/AJz4Mb6x2dXcwWD+0zAEc5NiGIn94PqT+pWastFiW1W9TVdzpvOx10dRWgYRWT7
wlq7X0QxY3iKIQ/Vjwr6j9vBPA0ZxomPIzj31UIfA8QxvkZbuCAEJjqE5x+1vWPN9ZNX/HfTBUHz
7iBEhKC5kLPdjTo0q6ucQ04qIfREaDQjbJCy136RqZihE39Ygi7WCZjfFImB4nyeeXPwVoreaM/h
AQU6W9xbxl9bAdgfDr1VY9rtXx6w9eInO4jCfY2g5t0rY+1umWwrBlLhkCHOTK8RvDiiThmr2Y31
zmN1+Ls4Xenw8FitfwdvUCPpZ39Z8p8Gj22gaVNBj0Kx9dr4LIlyr9Sf8cjTn85o+H/O0RsAKprp
gJuOUdQJseA82eJ0gI0BeFFcm+zIKJzXVkPzUH8vWOM/0J3dhhd56nIqjwB+arWd8AJiU5esA1wT
g+7OO+EVe5M3ACBP6aP8BeZXG7dcyM51L5SmyRebNI7hFJ7quCmaoobdz2PREokwLcLzfZffsvjX
NL9Bwcwo4REogMbRH16i63IQJBU+G4ZaLApq6l4gKgD3bBOwWCXc91XqBH7FzGUIAnTbZDUrtbj/
KL14m1LJ9/XxeKFwNXgznffVcNLk71Hwm/X0S85/kVRimwNN23OOjA4gtdc1OY61qjHI9XMImWT3
jbquvK2GkuSmHZMIHlOOxW6h4EM5P2NmVF4q+AX1bnGF3aPz5ZBumLiHzEuUI/LZ29jfiNQMbT40
6rMXrA0S8nljV+pTebCPQXpNBDdC2HkPGI+vRXiqJqvfID/l4WnDCg6lL9eGn1jXRvqDrp+cFm+w
L0Mlnsa/pTciuMh8wrteUXZVo8gSMsJwvjKasJ3La8JLPl5FumRb2+BwjBYaabN/jrsnfXN3gvHp
ZyroG4gr04mYEprc6AmqB7VQLAkWdtAsBmUt+mii4b9piCZcjNiifnkt+Ifk4QEzCjLchUd7Lp58
hQBK2v6ts5adN3QsXQ0AmBjzmzt3prleg/pLGiY8VvkTPyuwme3YJ1DoOpjHzhf7cR1NPGXrAg9E
KhO9wXPge6Ws73vDrhKXg9N0AX6fDMb2OxoYbJR53cXdfUBQx9lGTbCAYYVeTMSeIAn7cM/Wh0j0
AglRdVzHou6rvZO6F3BgQFyFMTMkMbOos6uReFfPxJyZ03AOYHshn/57gnTVgMTBz98sc9lyj9NA
/IM8oWWSGiXF6nhiVyUN8aelbA/bUETAugm6Jui+RR6X7JKrYrBSJVuKUmDE8bLd321nSNP+Xcm9
3T4y7jxsMwSn2Sx0JOKxWYVxYwlA8swW0EH6WoDrrLFzES8iGhPDlcCWmshqAx33RBBg3rqLMhwn
Ra4I1XTC/8eGpDFtcxL5QURNwD4nGmpVNYbAEnFQv7xqV2pG/s5nObVVIVAX0MWKbA9HsGiPAyX9
VpnJCW/V0RkhKQP4eljv47736Xyv4+zuKccsXzT/1YSt2gWMjFgYYNlNKN7UawLbBWwH4sbCsyif
cRSYNKlA8tl8k7mQTM0ijD4Rnza8DhxwYnKGhJClKaHWNRbUAjyG8+107cY+IGD1PsNc5WyCE3TO
+tnWy6of0Zf24Wdl79qB00w1QDzQIH9HprTW2YoXLdRgJEyqTHBONG9Y/V6ihVdNT00k9ZB2N58c
lJYIMfQ6fOT2w66LqMWubR47i3owollKsk4GYyH59/5WeDFmHMKkaIpHInQocttsSqYDK1puy1pt
sTc+b6zpaWmmyGTLkNHEC27lB2rBPHoFL7ictaunuPxpnkYVHuiRkfadBCOWzk3vBELOpl+mllws
66U0rJEdK7D65GnOnwHH7MbjMHLFESQYuDOvqASachOG+OR3OE+Bd6OUG09eYyXkjqMUkQeE/GD4
fv6QM4Ull505xfqeXXEpqR5wGV0UG4M0uhp5keI86Y3Bf2MxYBOMdMQohFU2z+rXhvUbZfY+FH5N
x3f/bFbggvBFBtn8GVDxGDpPIxHEtsZnZ9SYeNnIvWvV+/RoRafOQRslbSbybLgv8VgYt22cLBPE
tP2v7FQ1gZgMv9Jwjq/x/socm0941DZG+SbN0oM/VZhYn8dfOcTLn4ATmoWuE/gSu/PvSFNdSnwc
t8WV8bnhdIH6xXgz+xpDITmjSh2BRE7Cg84dwaopz9YeCofZUMnLm3+0HDLcM00IPu+BOFepNfYa
Df2pHzowrRJeRqRtIL1TmricUrZm71tduk3DejDaZCXpqRS7b4NoVHKhSfz0h49Zn7JNnIaTYZNF
U4mb1/YXFshoxFVBvmaqHPLnycPvNJsKP8lNQbShs1/orYYheLBV+/S+WJTPaaf4CjWvGwK3G5P7
cWF1aJFL8ODdLm94Hr6dYQKShgylduHNtJ05DvP+tKq9XXgr/LXSUD7NMylZWje4HwugtsKbPrCr
lZ12gBsCy6jeV8Nz/7q/EzqfxDNiWcBbqIJGWI9GYPqCs2eFAFbCLxdLd6nha9gpdTOrm1oTFnl9
0zl2L2bOKt8+zGhdvZ3tw4Xhw2OR7LqasAjA9/wdDvsC2tF+m9kEs+DlVTGIfMMMhfwewlkwWD9t
uVqL76TInlYNJdf/mur7L00th2Or+gEKyyl5jM3NBT2kMoqL1ZTyX97389OSJfDZAdiMr5W3PlY1
tSmgN/zv6YfXx/x0fRJIfO1Que5EWdLi6qvG0dZItwdFelZMNdJRXWPYTrUPCP0xjDWltcCNuQmy
3DI3dpOOYtPzFFt/4rZBGZT+mkV9UnHSwhSI9eInTS5chp0Wqpj2VuW0udYiwmEYFiv9+nGCvVz4
B4OuZMJJcXKPNKPN7vAmDDB4jUY8TrE/G9C6M5u4xZYZSI/kry9DMfaGyz9z7Wqf0i4VPJwJ1TIB
wjPwu44urwZDCIod2HJOXzA+V242hDA0LfWWMsTH8dMtKTYxIqKSQDTlazEUqQQMLbZ9Eddxzux3
Hk1Ic159XipazpJGFBYiH4cup8WpE+jER3jPzHppBlBZRkqQ6UO/9v1L4xAusoflIopI8isRpi8I
lxijsxVgrO1in2QraUBwU6Yqlu2tA7mVbT1Szt4YQWRK4L88Zln/Q4CtA1kIGB3nJ1WiCVAeb3MB
PEipBUwqI31EfD2cM8zxyyYY89OOkseeufKvdkvXjUtK/pEvzR68VOJipcD2HLJePVEG8uUssRno
xNhDYmg8hhfe/L5vWa1GZCBdx6imeC46TqgD03WnlLuymrN6lnxo+3kKGWlKWjqYqg39K00ISEa/
88Ew7oAIhlasKWnVvXZUuNGX4f8dQLzbuta+yUyPdiHS2TsIbQLezVymxbJwRc5B4DyZb9RUXMcX
SglaAAK6ESMvX4fDaavTmUyG2k31kWchdqNR10fWkccBW/nGcK4EsTLE3QIsqiMGQ4xfl2Ca9lfF
omhdhC0QEV7j1v91UT+mASFMHFn4rUeev4ESvT5kd025WWn1aWIT97SCApZwpPIVgjAB+VfN1MJ+
GC9AwXQXGolW1KpGZ5P37ZZ/TJVdGJh22RLPE1gpLvt3dJZ8cBn/OJfDjRN6hiIdR1Kz6qGr2zg7
j45Zv+vcXKXBLo+XSNkF8TWbUhmG85Mca2DvBS6Y6vnjziHmb04uyHsv0jAOmyIP/2rQ6wvxbKkd
OX5hhLeV/af8mm3lLorecC4fyPGaxJy68SLfFjWUU+lbfPmkBJ9mnb928PWtjPORAPA+99pvASy7
EtoDmEVL24a4OyEjePSVeFJsYUUyFT6vf0c+wIbP/vaK81HJUGa+D2/3rIQQ5DpmLGIXETks4DrB
GNFLhKAW8IB1qd832FioPDTQfrDkUXeWuUaqt+srChGEctXnsUdxlLD8wY9cnNFCBAT0NEvkpv56
09RZ4Y4l2kj99OhprnkJ30lStvYNjt5nDsuLa2KhJ4fSMYJK50n1cMEydUNWljUuMjLwfjkfvFrF
tBgUqKn2a9682S4OjquSFFLqWufscA+cFhqsBx8XpliE8KeXG7ITXkk+aO9KcuLgxTc+cfQ3P1fY
80gGKmtc1Rb4RHrxxz8fMyVuid+fOZpyVJVGlbZzMYeCVQ7SDbboromaurNGTNM4Mr8vLRaJKls9
VJiETAREL3Wzk+gi5wr8ekQlKwO7ADqZFFj66ZfTRrsRKh7cz7/MEt9+uI87WkJZUygAKCLR9t0a
xnU6YUpIOj5m8rcLLRixogtj7IOYg6n3/1Aw243np16AfNcvSsDR5HiCe9osq6Rdh+zsYsmH0YRZ
3tjMFoUEt5tyW4UBOOBxnGz4O9kHTAZQWrta/J/ZQ/QS9+QBb93gah9mRmZXNFL1cBJSeSJEZ7aC
nBQP0hvjgBGmod4G3/JHT/aWGLfyWK3B0VoPAMuJJuIGJLXjDiKOGo7IBzaG7NQwC3O7GzNF1SWB
yDA9qvBts/AgC27BpCDuh+w5kyRM6Hb99o0z8FZB5Mo5I+P82KdazJTxjwm9KsV0hkYcUUggOKef
t/4EugrL+/9WS04ZL3T+JGnH6bCCkQYfXc8ETeN0zYW9IG25zIZctRmfgkzgFBLx/YfB1Jl1GRfK
3+ACAxll3EOX4OfX+GNLWe/lDmfuf1VK4EmgdpHgjO3CeP6GS8mCBbesvHe1nFE/t1lm9pg1W5JJ
BYMdiV+ZGY+tWH6YSyDZ0z/KNSZ0FWV68XoGj+QkTfV5QV3hR60iIMxemnowtgciW/Q9rCT0fEcJ
6S7prF7DvDci536fgq3r1Jm8drjEjJL1zm3DGieu2Rtto7GfjQInv9l0oPNpH4ZKloFAi9rPniq/
22qdhTohdMKbl+TjAxPBuwXpEHQTftLUvHfUr0EWEav/Z63TCI8K/tTvvfINBMIzHlchg59zyfSV
HiKe4sFnfADCRiCfW0taSOJ5lKNEnBDfjgd/0x1pCgYOh4Jc1EF2dStB+wuJHycjyrvXxGJHYZey
CZCDq5zHrgajK4/zkmTTZpIByN9Sk3omsZS5MKKjCkdisvNjAwtM4aYiU9ZrJWjCMXZUoYjVtdYz
NwOrTpCg+hr/XcCbl9ypavyVmRYRzhyIaJVry/ON7YecTZI2FjCJhPdI69to2NWqNlkriYTaatB4
Ct3hFoiaERcQcN7StBPNpL21Fe2RxrAsf4UdFbVdwjYpYGrcQl1Jp0f57OuzeLfXkUGoHA+8Q8Fc
1boIj2JwvPEslslZNObwq1Cs0RqdPfmm9eu7zmaBdayP+UJ9Ohh22yfGePGozHsDeFd3dfaUwMFI
triHHoeIeidUmHHLjryKyohnJ8esJp85WjuehIdjOsgHEb3s1C5MbEZZdqbV5gI1w6yNstK2LC78
vFda99nSW6bRu9GnbdDpWEvurrrXAHZKMGavQ4oUeKiNDH2wbVziBM2PnJEwVMv8Zj8qnS0PyzvX
hYVnBZ7dzxbAo/I9DERde1+ls+hL2KlEQ3fvioeUpBL3Z5i9ZXZf5FnTPEDjhwDDftwqasyLveox
OJmJWmZlwtlkJqJhRAYqHNoZVZqvDLRx034D4fJlYy+mqPB38+Gt2grO2d2pY6RN1Gx629LCDPQ/
1gY6RfwQVbyUAzwgn3Z74Sw9zJXAuw8MJowkZ4+hqicLI3b0yHZNtG6BFX1gQ6zBvfpnGODQ6P6C
Z85iVjtkjNO20xqiIbeX+LAFiwDIMpIbC+txuv1EYdoqI06mSxuoE/2KVEMcN/MAaoO2oS6X7s/r
zxpRTFyhgyrsi7D+zyC7r5Nf/LHBnQVfgDgCF57399vCj/hNkV5Rqf2CW0JQcHAU6pxPQ414aZ+E
STPLQhfcgtn4GEL9GIT1hpZhBjmUjt4raXNFWuxbx65ORZJKFQApEcJZTVyNHplKNcDQdm7cX+en
Acyggzevp8JNn1OfPvT007+FRlUaA2r1UwlkZnw6jEXEkmnQLPmZdCRRdel4vgXYsTH8k7LNWHBJ
0ummQ5ntKLci3O+dCS65lnom/+WFhTBKBoh4zbQAXXYoYyQ5eTvjufKQsFD4spOjJKsZkl5hW8cA
rBgU/fcSMFiOiELPQYfpJkDVEHsL/urP77EBHf0jaPNlM5XtZ2fRSgWqiD8fXtfO0HHVRsQ8fnce
FuUF0thlvVJQVdtmPqYlFFtWho+stQw/3bqFXAX8phGCqSuz3bbaWoQB6DbS5t3Ulz+5R3jCPdEa
1HDtWISnE+TLbbixCStH8KExmrwXtUsph9fLl9kyZdtYC8uGgBsz1Swg1bFbHhHkRFoXQDX7Brjj
3tXQeTd3oVshfOhFPeRZ2pKC4Poot307arYmiNAgyoV/NGEXGZ9e6D0hgWs6Z2c8KwoavMaR9iBr
NLRzg52ZA0u5n+H9JIXPoOG4f0Onw3OoQMm76tjeaQWL8i7poVFb1eREj7xZ97I3JoTftL4PiNH/
e2UdyKWGfYbun67MqGTpxQQpEdZl3GSVwfEmVTfhen5ElW0u3pjcyOgDwkbjC4WzVTNUdLEUqoii
3TTwpllrqSUxhQ+jiID0bi3VS+mfFNKb7DyxsOE8/kKyzcJxDBIAmGzxXajNVagLLXKt9/jcifxk
cIdPc7S6/hKsqul80hbVqFQlTp0zwro/3VQuEra30F5y2t+5HHCun2QFK0P1yIDDlyS9BQ582zlK
qSAI+vQIzW9TX6WLH2udcW52MIcI/KFUeC1fZx6oYX/Hg426ZWz1OGiHbUevW92TDA4C7xvR+7Xw
8w9n7N1GPofHcyz/x3vFXpX6HWvrLVtBbqWVhUuIdmoIAYmjQ+walr8WYMmN3HJORBmB1+nTqUSH
DmtIEYoyaDrS20mFvD2tkVNdKl5+UDeARbxgoF8Hn0dlXMbcAzfSF6zwhgt60KAefuXKbOO6/h5p
Nuv6syn7TIpAUsiXVIbaYMgrQgfWUcNxZGc6FuerXPcnJTW8g8Uht4EZQw0Mg7bs7IIIAjUyfnfY
o+qPmjtKjYi1DG0QogsyP8pfrK1hIL3GMkEja4G9Tk0SLvaP/Mf49UvcSL581nNTfnfjmCHw9Ys/
dMGbgaigc/duPPeGDyP8RYs4Z3R+U2YT72Bh0zU0RDMQGUHZE/8jGjJBd11Gx0xd5VqPalBcuAOe
ImMARhMiWbyfbidy6Joxz/dDkYNzlO2urrSZyaVn+o6o7kYJpCwKbGhiGiVPD6ofcUe6KJFI7mDJ
xuP+gSyvD3K09gdzbX0rg+JeBCRqOAzn1npKxHwuXTqz/wkdQRAetDdFGyMF9mb0WBnfu5Q+Zy8W
dVXsAoPD675ohqDKDfUGRE5tnOqJfNXo0DQbUVWuJdnzlt/IfyDlGXnGBhodXMIwFykm2+xcmNEW
puYs0bkcv0Pt1QOSA53SU2oXCe/0hjUp86ZKlztFF4WR51B3rD1+slsCQcqgGM2u+xwJxH92T/+C
LJ0EEzacRteWXOB642p4IEWjzUQtqB1odpdhkX6nI5zrou2zfMrvcpHlxNjani5Pu/EaGx6CDJSQ
V4KkCbyZmNaBU/ATMIlZWnY2lh/nm2SgdYj8bnlS3JqLte5imDXgEzSM5xO0qGH9CniLWOejnibq
ydBAiOXkHx4Cvgm+m8z8TIjRxK8FUfLCpFYKO3O9R2J8MGt3eH9xyQDXYTLX7D0AigM17hk4OEsT
eEhjD6XreAJ2oGb24PgqxNQEZzdK/GQuhkBMRgT9Oyse9k3t/O6gwWYNifm944OBQRvZxl9LnAry
M0d4z6toM9x3IkxPuObw0q0J/RXTv1YHy8FTkddhm7ZX03I53Srz+e6vzScO+CAOs6t+s1LdaEe4
Tb80vb2LYT41gfb0rgbn15exGxDhoFmxTAhWqmmTj8jmxPk/NdWpdZbDBLHbB7IOdCptiNJOwy4S
xvhq8sOtdmjry4QDbdH9z5P3Xb6kIgM+stsGuqpdtwqoE32vosnzQcfBygnL4hvba1xo1FvcQ8Fg
XxwSXhseXse+oxhxqBJLp7lCLo0asgP99f2qznsVk5QjBewqaDA/AFOpbV0uZQsDyzs/SfLUgoAs
pgBxKWiqBp/pfrNNXdfV9jTfyRlfOqVAKFaBUIAZwK0mdFH0fbKeOanL7Yyovx57vaqvhtBjj6VD
wuGiQxCqTJ2Q+4WfxdaOc+I2o+cpk27tWa6Ga4z6QInd0DkejDMe3NcyjHYUKsZhnPILgYxtyNPI
NVmSnM1gGEqyg5UIToLUy+eCup9R5v0Sso2J79o2tsu8dc5DkFQxuhDfMAvNBY+TjPiPT0pxKVmA
XjyD7zN83M8wQxdpGm/ePCANN9XBbumGCTY6O9v2fkaRWt8SXIYWWEavn2Wl5WCEM6TQGm2jHPKf
+OSRbqQloBzNAmT9uaG74LtpQvYO8yq5+Cf7O2ph0zxGnEdFIt9WUvQKi2o6RsxQ95qtO+0UQVIQ
MHc8bFoZs7aM6HD6CNRilQ6ie9zX7gDll64BGAim8nO8sm7G5dqB5u/k2uRm2rASMFSxl2xT/OSv
Ga7NjKr8y0Rt5T+6UYe39EL6ns9wTb4jz+F0n9O7cqBtHHgCT+Jn60c/s0t8HEidusOKQAQQTsWx
MYBEHwIEqPKHCxq9fLYlb+UanqtBmD9erqf4vHpL26GXDgz162qmO27ilR9xrUiMZEwIA6NPIlOK
FiZeg/qsa2Vx1Cwjnf99E+I7PILZvyH/OuJZxCejViCHKs74GpgKXF6SHl94z8D4LLLuSVdGKxqi
MHQQ5tx88oUTtKeNX+ZzKjW7FeK3BjqhDJpervLaY6r5hUtur6shkhQYXESCD/FWfqytZrqUbECR
y6CVLOrb/PUvlHK5o5yDexdWoZZtYaU3A8nPF91relXwDxGaarJ+18dXfbOaCtHn1dVlaA/RbMFV
xo3bXSHfUTHDn0VMC/HwAOe5C5z72gVbRG7fIXQQRM/C/h42MrK5T0y0jDru+a3ndvRE9Lv8klsa
fpiJuMveCLlAxLdE84rsAFbqit6eslxjqwoZ0MO6fl9nY8omwoyVbwbfAy9e5NomJA/c5oggE/0O
LL9uw/SdfAZSRa+gYKCzam6z2Oo8gzaHbo1LE/FAOpTf4nttNVGLAwj49+YbbjYLnnmQUrpO1a4k
7y99WY4BLHH4Llz3dUYv/4bcBlSqrBLqyJM+HU7WyNH7o9MaJ4JorfxTOQf0Eu0D8fNkKp9Pwul9
cRopxpGVxSjtAaLr8d9Ok32073rtQ188UhCQ9Wc+vk81kayHLabruUal5a+wPuKd1TUgH7q2H8la
eGO6Ny+bTKquzdhuDLbl9TpxfKPxjyh8dZX/iZCYe5S9hC1sjv1PNni9j5z+oropQJ6D+lbnZheR
aAv3isdcZK3mgr2cp5p9ugCw8HYkApoLvS5Pi3E5sDbQZWILk1RxdAJF1habiVeeN7IVyBhET2s5
C46aebgHtTqy/h6F5jpIxQBFDJCi7c4ZmppZsX/Y21Scg+1sf8IaCuk3xDVQdhqJAj+IEWQfZeTQ
quW+PZmU43HH3874lidyrJx9tWXdIDuvD2L0AUidRulnOl98TkrtjFDFO87AC4DhNsmlkizB02ZQ
LVNnSoJhQo/RDEzpFbt80LOnpqi8oLe5EFn2EACIfXLSbA/y2MOXJBqDxgswiqcldEUKVee1i9pU
KXxKktATtKj4s96MCuyGUYrfkKFiFBDaNAqopkTWc7YfYFzwx9BwzfX12gmrJRvHrNd/Usz5hJ8K
qEc1TqSftybkTEhIndy8r7spvri88cEgaO3vxeyWRaWrPtXbqT05ugiwqAUN9bwxB8XhJZqnnzn9
5pZM+58kGqi+CUC7jI565kl/wrC1Dg4yFqtctk0TnJ1EfzPH7KRMzZwfoJt2GgzGxeX5KgrjoYGA
kiQLYvQM92WMWWX2xOGgUL70/BvZbeKBtjt8psahS+piFeoCZGpTg9wXRgpPmjrlfLIF3h1FSA/A
J3TOwAHdcKIYEAxZfEtZE+mDA68uYJN/c4Ru+NuAYS1VE7N6gmsnVeC0Ne0DVT93pyE2x7q76CpN
NtK3LHYqCPoK4Fr9dYyBqVftT7KDaoq8DQ9dw04RUdfGQfl5s5Y382sitLCUlk67uiDvn9MqUOle
ipKr7iUFLulTxo6BMNx9/tsbqK2uZPRQ0ek7KkX4Onv5ZWLGhMfMOU8U8ZgHKLaXaSCTwj+FaVXC
m0h9cyTviaL5ZgIYN6ZTtC2LDAdRU2mAbvjagENb++NDdHsKaiUarP0l/3t3+g970zk4fNJHJyHr
pUbzwLIL2hYSkYMv+ghB+ghWcRbF3L+GVC8Zd7Cosz7y73mkZ6Y7EY6FCVEfwrmhWL15QNS4JKEM
/ubjtx7h2Ibd4ZtE0L8uGj31npxDtuSyQLDeA7ogHip3fDCBrzepPKVLgGpu699twMLiNRfEKirV
owlfH1Xf191zcTaeGndcI45MOYzyH4cfX6/xtXZIZC17eb8Tut7EMenRQEvOWWPv/KVmz5Iv0VBF
rIVYGL8DC8W37nFsp9yiTxCNyV8n0GMXtmfx73O0P2c8oSLGf62h768K4WOD7BnPGSeUSVgKT/MH
20kyHS+VtTAhoHfBQkNoCMJ5dJeSQ5w12YeVvxHG9bD4xfZMuQ4ckCfgm/SIipHNXUuZRSMcEAFi
c4SshsQk6jR8uvVfdFSGTBfSubzfq0QguhbRT9uDHWgQcD72mAlEzkUO2Mp5+08eoc6Uiuce3Q+u
fMkUtyQXZNQ2t8e6nkt2vLD3+a6FZRSy05OTKweQBWaKXkI8B9fddO7xKoz+BEmDC32sNQQM32Ud
tXHH7zJ+5iKzKCSq5rGLdOZ1/6eo4g2qSC56G/gEjCalbF1YumhBQOyP/Q8iQrYAa8oNQ8kpIDmu
SDBR/zT0v6MzsNGVPeTJ8IZ37+awq2KvhLcI56nLphcn2TFzr8uWP2BGjY3l9daf8yA/8n8zjMaG
ZjxSzhb7zuBKgTmKJJsQcBDdPxqPBcMU4ne7xnAVyIH2pLUtZ5su6GH8HZouMhhI1u/fVbaZLc6N
7GfSXGgeuKFxfncBRoEKy+D4G5rBVxJhvxid5trQ68Vkk8lefVg+X7/APqOTq0Ee2Vq9DdtHhaeR
c0oBkqF8ikEHLYXz98ywaYjVMmisCOZg7KnSJdKGtYxxliRn8ZO45Qk7nxJfEu10sDm8h68OM6Ro
kdkCArv7stvxIZEWXhDE0nX5VQ+Nb8BW79jv/R9kO9BewDV+Y/I8f6uCP0krS2+gOqstqAIQPqT0
nWzobc4eQ3Ag0zaZ7YUgIVH/hVeyngLT/pnKzq4l8nm5FsJNnW/0CEAcH3Afl3J6Dp+S9cH7+EZv
gEHUbdbcFyCmHOLl1NB9xdcvWHPYvLcodSyHV3L9Q7B3UEljGiKvNEYNeBWnNv/zX9rPkLv+OOM4
J915OaExtgVFIlFXZsGumsQ9A6mP731T94fn4ERyfFneHP5DueVVoMvE7poqu9VBIt10gIkmbzf7
skuCOYTX5BAU5IjJe6Kq6lGywo8TFdDLjbSc9p6gw4YYCm1qfFbCiOUscSWj5jNPJa0KajrEZgSQ
ZeSkZ5N+rga5Ypo7BM0X9eRcbwo+xyM18+n/DoIHx8lYe3Kqpt+XaHk8bMf+LsX4ECvD7bF25RRD
WfXj+DSSfIKBy/k4zTnK6B23ONH8G2YvmyRYnd+ZkjUBw1g4nIjitfLphlL4uu+7GQVI5p2QpneB
QHbE+wyaphdF82ZzymH4BPoCY1sVaAFKhKDBkdoHIyABT1n8KuFHOjd5Vc+PGyXztpbdTB75ZYCp
my/S5BJ7lv3ZUlAWTMsxciKku1lKD9HZWhd/UHZWGfhbXkRp1BonKARwM+W1Pf7Xw1aQtg8x1Cdx
k8i3m83OXR6qKuSXvnAhb0F9SYAWs3E02awwumOdyqk5x5zN1cq+2W+ClNN/yNqBrmVeeuT1DuQC
7ZNlI4HQTBDBQl6Mcbk5cyI2Yr9j2Sq5yzgWsXvLUyOHCQP+zC1CcXF58sG7eahscZG8vUVhTfDU
RB9VB3f5cUvsvTkcCr633Kku65eRftIDOyiOO9CiZZH2W6RNmqk+FDRnnv03ykK0gpgH9ycIYs1X
nKhvSTfILaHpUL6vByp+TDJ17UzBdp9ZEBV93GPegZAoYat5oqG3C1AZiVkN2nYKdaLeq3i0Viz7
Bf3YTsc6QFx0JlH//C5NsiNgeRn5rTZ0UlNXJMUVxVwcTQ08XVfxpfb0C2uNfQOT2bCRco+ZwbPd
Qj5CQP4CbYDw2Icg2JjNRbHQxrqQ/ZwAhIK/3vqlIxLD3V1cJnZQVp01zJusS7J320h4ZUBOy/Va
UAFrur2A7trt6J5Vh6w+nRGS2FhEIMZuB5RDXtkaQDBxQUf/XQoewNZwTXb5DzssFPACdUPXSSqH
DQohWiXyDPUVVowMwnkOMKOEueNiAiMqxUesv/tr43GMO0q0CQpXaDApBE/FDxW36hg6P0j/fWsW
XRDXp28i6Ajp300LF52iNkI2RC2Mz0XeGV1WyxoBZGPD9GRgbUe4fQq1ZThTp7YoOn5tHTiVHdmH
Lh7cUHqH0xdQy5pglYhRYHF+q1WzM/xu2Wf5XQWHQZlM/QJPBTV4wkY4u9D5iJP96OZbrn79z48w
dCPuBYefJE3US2rV6IML6Z50J4GjrRKhbIF8pzqFwgzihSwVQDZaBtqsqGPxyWQ4Yp6wY8gbTBwd
0e+ExGw+5mgM+TfDwctTk5Pgr3BAVEpohtR1lHlbLXdKarMfrwtBX886j+80eJStsGPMcMzMT2yU
7EUcB/1hG/569jlGJ+WzcCIMpTirj6uhkPrKBrxt34lMUrmxjSYeDmxRvYlyfM3GSPRd5APDktl7
YvMdGrVwq0On5p/sxLzGMtoIjOb/TOEkmx7yTz2jPJDLdes8xJMpGjjxDBbyGHhKyxeb7ZWZPkPe
YLoDyCLLz6ETQyz3EiIgj4EF6kAAHZvy/qDKC2LalfUjw0IxJBudo+bQnSAQW4v+UFfAy6pE6/TE
pr5/xCi97VopcNjKyTjBcMa2SAeDGnZhho9tVLmcx/D62OqYZVi5lwrmDLltVLBRwqpnJnqx8PXa
YwBMN399Kpzkr1UNUisWQ8WWuVXKZu4Gn7CF7/JRha5ZTZdfG2+1ClXNezeb8f1eJBtWbQBiq+wn
oIRamQHCAJGmVH6jdQqaWBD/lnsP639apx0+6BfvPbqAX5iMO4K0KC1tbz/sxfYvAzWtCYFdAcae
hI8lI9bhSdSN5D0HOvoyI3ItTQO87CD34Faax1xy6OhXq1f7dercvjliIBqF0CcktxQGXYPm9Cdv
VSLg/el1nBIwuAPMaoh1SdNDPQUQX1Q+FTIUliHGvBzayNrIWqLtSNJvO07042hikCW0uEhL2QKa
6uuyne+g+TZb4qInqbRhLJ3z322w2bLNbs1mJPOhyKCLpMASDdWem+PKhq63My12TRS2DYRtdyPd
LquhPf0rvMcaLp2g1w2Tynql5897hTesQmLGT3dMfrsyVfDNxPT50xLQOHAzHQZ0wPZGRQ55bWZX
fZCZN1h/kWiMdt9DAZDaSqoAN9mYBwPhs9VOjeQWW3oF1d6s+ZZpr1liZ2zzNaxXdqo2gvjCCT+K
rj0+9wFkSX/l+u0JbfOYGRgC8aXrWZl/Ihf+wlU44R/mIFXjudvTicZ7u+AVxNmMed2J6+bPdltI
scDPcyY8Dv6n9UGzbnS1XSFsq0z0y7AaddgTnJkHTvySuh313MpnSSQOzSggUhFvUN75xXrCB/UY
dmre7+ta+MWMn9u6b1lk+s7XMUR0PoLGGrU2KfkdJLZj3OUprjSFxQBJpDQKiBOFEUvU5yYw8Rwh
2lUIoaxO6CBOEb9VF0KPeyKAK6uMlhRFOlMxQcoG+OxuvaMKpLHYOo5warHgrfKMD4xFyqdtv7YM
QQLa+6EdTvU8vmAOlyNntP7BD+1+ik8kcm78X4g97h296CTDHuV8MGWEDqoOkM3e+12+6VeHhE4c
FRhpUHNSyMD7nVbVYFRMzd+RqaWSlz8e5vaodSoDvCKK4GdLcyjr9BdlL3XX4x6lfXn2fcpboyvF
qcfWWKTKpuobFqBAiTmweLtXqkzT361bRjNzt10ycOhu3mqywnSZqaQoRv4jgvLkOxBE11qZtGsR
B4khw+mB8YZkAj42FD2rS1XXxj0CttY8QfkJaBoEEvaWLmLFYzFm6ux6RPJ4LEbWdgDroNh7t5uh
1PANzgRc4jjeCM0hH2Y63puOhf+FTs4nmHQQrMD8F5iqTxlqYtaF8pvD1P0S6bUN1o4X0BxTAgpE
uwVEdpNgLdtnqaSsZ+fRPTeqJ3Y8rRN6bCALOqzzs45Kx44aWUSNqneojprNV497sMBciu0CMD8H
FocJHB0kPRaMBoImcCu9fhuX3oM57YjOjZEuRIwBaeNcVIHrYlgDfEKALZs5iB5xloUDEV7IYq0Q
ojuBWznhfpOswEMXclSfWgEIGgNKY0dvLoj4zPEt53Y3SZMVrZeIge54SQxMQUQsOzatBVJl8GGn
tUr1pxcVgpcqXrqFcgxSqxL2r0vDAc3593cuVvytltWO9VqU4wBxJjvdDKcfgZ2P2+OFzW3g9hbg
aEA9OANKsIwgf+IBlV4SPnwvlvsFt1wqjAQbgV+EXSJT21ZYKHLpIQD5pqoZC2HCt+JHFnZN7Nki
b0L1Cv06zpUPpZs6zBkhns4m8pFqgwbq1DHvBS/ZHegaNEIEku5B1sVPDuVyn8xkY7nZjOr9rGSW
JF7gVPG/8ZCa24J6ZLxGPlpkclesjpnxhHqm3ZdCrKobTQMQfQxQ7crJuqBRZJfU6qJfEjFQIPRn
QukQOacWwpQAmnP7gyuS1U63SJuq2ENDanNVSZPLGmNcOUyUCyLgcE5mYeSgTqxZi2kHWnc5DiCI
cHDL7OXUnFtJmj0cQjdi3gQUUZLJxmgn+t9pR1vHMrm8RPTJrRh6YhJJuKQU8Ya7+lyW0qu6waGt
PSOzTYxLL8wFodbNxXYXFJvvz+YApyIlAbGPX2n0CQp5UUORXQlVDXyD2nAEYuuuEh6ty/5V+0Vz
BWHGCrF5ScpmtFXnNAitgS1r1PqpdC+bZAbm8rFA1kBZSE9/xNcnCYWBoYC6TXEx+84jDU4FQk9a
9+XMaT+Al9uEeNV2Oec7fE9G0fpSSVjwffGP4GpiIr+LVrj50EXf8iHopdC1V9yAOcqUFsUqQMUA
n6nmxSj+mAB4ChmdBWWlxo6MN48s6k1N6w+yJQE2zuIunksivt+uG/9FxxX0VRu3TRGexS/Ba3+c
hzc+kB7Ny/m94GGG+6XZd9rnEgvr7TpncT+/xxQFlU+igjlH2C9IO9MEW8vnm1CliYvq2HDFVbC4
WfNWODcatYs8SvRQGdUswV7X4MZKSw17CyGu8gUBoLZUmeGF310JKn0q6UAlFW6uUvyetwfSInG+
JjiWiW/K0xm9iELA36FYS2vIIUTRBRC1TuOWq7JFbTBpRsuLF0LGp30Zv/OW2RCC/n+XPVNi8n6e
USSUbYhieBrK3m8JJF2k8eV46nh9UNS2w/M/+TfEqiHDnONvvzLUjMlejKvN93CdmCJaYs3HAkX4
+E83ymj+6jkuxdC7HK3xeyzGiqdC/6B8yceOA3GWtdaOIVWlloHBaBgqoOVu+toPKEUaFGbrTd6g
dh5VJHCxAD4SusdDwDAdmvHJ2ohqjnzVDVWG9fhPoy/nBMn/6SeM3QtXhUsyYgPwuvXx+zBMTAmZ
qoanDoumZ04iuN6sTLG0i1UYM3zVp+h3FE4RGGB+K+wuJt866ukYDyELaqxWVZ3Pro6hcb1BWNo5
5DlmcYfvACJNYwLHYh7Noq7Cnn8Ylddu89ZF5mzouEgmZa2XLMvFAeZCs+sd9mFDtpe0TnlBqIhb
zNH23w3nqQsXgjP2xzyZdKGfNxOGrbm1rWsZ/e/OBrXnZdW2tvCpBTPDSv9sFGgm4Y3wZjg+FRa7
xitmvEVZmuw5m58vr3UK3NYKH4A6tfOu9NDdbKykPEeEvtibIn+q/q6WU/1gBfS+tjxUn2k3UKBp
fh437H/AR/yGvLpcDjq/nYVp8iVn+baKajVlKboU8148mQ3+NVxc1dqHpl99iaEskNQvFZ/NxH6n
QrYZDYgYlgRCqXy+8+wJ/Zh1LZ0y7BqX5sdoqqDTjuoaPNg3YONbh3OcS+78ocxRJoxNgIHGz9P2
4yHypeuqXyWWCP2AT9nNKUhhIJwXq4eN2rvqilsVyyFooNXPJs+2CbAmEFstGVSQ2yZ4zWVJuOsF
ILyJgU8yMJK+79sMmML4BylIXh3SQmZzK96ZMFq5rWi5yquV1P5xPlBMM6K1gmG/c5MHK/fx6hwv
Qc/ccNoi0e5MV299IMEmE8smFrm0/SV1GpRCf71MtrmvoUlEJYS8RQep8JBm457EW183KnxJygE+
UjTPAZOENIsy/doKamJSsS4mKTaKb3vwLlm9rXxX8IEbDNN18ganWvinkwCDk4fI8f6MJTHmAWu5
Rz7/hPvbf8sLqaukqYdEgqbe3AOu66uYgijLylJcY//4EgiwLH6aRl6X1ZtWasXkxI/2wINqwzIp
Gv33JiuzWWVMYzb05FVehtiG5BnBrogmyTEbE5nms5YkaL6i2auKa13np2jQHvAoxxjf7bhlgjhZ
C0mT6hSOlixMqX78f2GHUCrZ8n7eFCmaSLi8kFy/svTcRvO63tq8cRJ4qoTrUUc14H/xtUZV7+iX
mj2jBEVfkXJ6GQ7mNMvEd2kOOhMmvTPi4Ol0ruf1RLvpBfl7biQjGrxdWYYAzgS4Hf2lmnrqjpZ1
CkL1Wycpddd7EMr30iH6HA+Jx9ipqNtx8c+xgJEy34zddefzyQsDn0j6rLIDSfpilY4q/hFY9nps
1a9VKbKl1y2HqR9HCRybac87mATPAPLY4ramWGydvaWwveIcmK2lpj9/emBRbsXvnetu4ja91+nj
c07RHOv7q2o6J+e9J4AH7Nsdbr6LRRY4KmpGIrjxpO1ackzaK9F/dfvkZhlwf1wGS0hl4kSFJ6CP
PpHqS1PNSR9a8e0Tn92bf+HsqNbIUhygkX4v5vu5Fh2ZygKGror6FPp9i97eWf8H7WXxjoQDcxtM
M/OyvSWlBPlsiGMN9x2hvWzI65ehVTxlpwqKlTy0axIPRPboX9jh1kHBUROCraTg3wVENpBRqsAS
EZHmaEzlm2YJnkdlV9rlZ+AQl7H8uS530l5ijF2hRRr1onzKT7vUwmkyBI5xwx71SfqovEuSlM7s
GXsnMEY9Ov9cP9MvWZPRZ+P2TcWFJS5bKZ481MMhmRwSjjqgDlhb8MlCuMCYb8xnoTcnDApVGQiA
qw3AiXX4ON2g35gtnpt+Hqr6iSecTPS4dsHA8ay4ya+MyfUOzb8woN5Hp98lhctbAoL69boyJpLH
A1pMKsvDUil0VaVq4e6zgkcKhW3ILfgFSCBJN6szC/fXdwqk5qX/vNtrb0LV5aUrVFbs/dB2trQv
J1YeFa/C/sT54Bfa+bHhRMvb6CEFo/MxZl1Cr8+x01jiHG3KwcoY4E6JyYKGLMxYBGNtPYUp+yVo
TWZbTQwnrTPlwFRs28vAbp4lY/ngDBQJoAeBBJO/+yFQJfyH7dZTnTbx2oVqlR128bmVKh4mA6aC
LdtvMUaipArw60SF2ewL+MgPzPntJblvciG1NbMH+ksOYouLq3NbcBlJw81PpVWU56+0cA51PzNn
xn6JDX9dnUHZHhj1cfH3E/KmX0spaZSLf946R3RiR0F+2wYzEn2YzhfcBi5ljD0wLPxXzxc4m9Zr
R+3N7tx08fe1s+DNSZ0Y3cCFl5/nGK3/V04jEPCcb8QR1cHMt7Sf53SiEWctdv4JsqV/tytq02dF
9fkgwJIG9IMIIp/s4jlfNyUGoOZ6Au6AMz+X2zoToKcu9IatovTBfvkxx4P+R+j6eJsobmaunEGp
oegBHNLlMPpQrz4j7hZ7AOvRhQJZLmSwNI6wzQX7C7tAezyusw64AwmTUiz7PNvNfISshf1tTSbM
apApuIAFYzyGWRHqNpaUnGoTvMnYuZEOoZYl+04Zcw4pp3nfckgIZJMq4glkLUgBd0vsPim0itod
M0wudMdKF6bmWUesFYcwHtmSp4XuHbZ7W65h9hxKjMe2ihpfyqx9SpcVm87LYtUGAgo/dIB+DecM
37pKioCatDROE++4pWAkyByaOXVzazhzPw73djlEqcfqGDF37g9udqHopsrIEV9GKdmRt2vMjj/L
DZeD7g1BFDmwPmaD+L+vo4V1X9Sx94NfyM5VdZ6Dg702TF3k00JyaF+jV5RQXGSZajE5gTWySIUn
gHZYS5muHq08ivXJvKNAzzzn9sdLj9bt+iMJo43FWdOdFsKfllIdKMgCKadcqgsndcK0FKz7wSux
gYwteId7Sa/t8NggQvpNpTU8lL22MlT2XA==
`pragma protect end_protected

