-- GENERATED WITH MATLAB...

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package DDS_constants_pkg is 


constant W_COS : integer := 16; -- bit-width of the LUT elements 
constant N_COS : integer := 12; -- number of LUT elements 2^N_COS 
type type_a4096x16_std is array (0 to 4095) of std_logic_vector(15 downto 0); 

constant COS_LUT : type_a4096x16_std := (  -- s[16 15] 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111111", 
	 "0111111111111110", 
	 "0111111111111110", 
	 "0111111111111110", 
	 "0111111111111110", 
	 "0111111111111110", 
	 "0111111111111110", 
	 "0111111111111110", 
	 "0111111111111110", 
	 "0111111111111101", 
	 "0111111111111101", 
	 "0111111111111101", 
	 "0111111111111101", 
	 "0111111111111101", 
	 "0111111111111101", 
	 "0111111111111100", 
	 "0111111111111100", 
	 "0111111111111100", 
	 "0111111111111100", 
	 "0111111111111100", 
	 "0111111111111011", 
	 "0111111111111011", 
	 "0111111111111011", 
	 "0111111111111011", 
	 "0111111111111010", 
	 "0111111111111010", 
	 "0111111111111010", 
	 "0111111111111010", 
	 "0111111111111001", 
	 "0111111111111001", 
	 "0111111111111001", 
	 "0111111111111001", 
	 "0111111111111000", 
	 "0111111111111000", 
	 "0111111111111000", 
	 "0111111111111000", 
	 "0111111111110111", 
	 "0111111111110111", 
	 "0111111111110111", 
	 "0111111111110110", 
	 "0111111111110110", 
	 "0111111111110110", 
	 "0111111111110110", 
	 "0111111111110101", 
	 "0111111111110101", 
	 "0111111111110101", 
	 "0111111111110100", 
	 "0111111111110100", 
	 "0111111111110100", 
	 "0111111111110011", 
	 "0111111111110011", 
	 "0111111111110010", 
	 "0111111111110010", 
	 "0111111111110010", 
	 "0111111111110001", 
	 "0111111111110001", 
	 "0111111111110001", 
	 "0111111111110000", 
	 "0111111111110000", 
	 "0111111111101111", 
	 "0111111111101111", 
	 "0111111111101111", 
	 "0111111111101110", 
	 "0111111111101110", 
	 "0111111111101101", 
	 "0111111111101101", 
	 "0111111111101100", 
	 "0111111111101100", 
	 "0111111111101100", 
	 "0111111111101011", 
	 "0111111111101011", 
	 "0111111111101010", 
	 "0111111111101010", 
	 "0111111111101001", 
	 "0111111111101001", 
	 "0111111111101000", 
	 "0111111111101000", 
	 "0111111111100111", 
	 "0111111111100111", 
	 "0111111111100110", 
	 "0111111111100110", 
	 "0111111111100101", 
	 "0111111111100101", 
	 "0111111111100100", 
	 "0111111111100100", 
	 "0111111111100011", 
	 "0111111111100011", 
	 "0111111111100010", 
	 "0111111111100010", 
	 "0111111111100001", 
	 "0111111111100001", 
	 "0111111111100000", 
	 "0111111111100000", 
	 "0111111111011111", 
	 "0111111111011110", 
	 "0111111111011110", 
	 "0111111111011101", 
	 "0111111111011101", 
	 "0111111111011100", 
	 "0111111111011100", 
	 "0111111111011011", 
	 "0111111111011010", 
	 "0111111111011010", 
	 "0111111111011001", 
	 "0111111111011001", 
	 "0111111111011000", 
	 "0111111111010111", 
	 "0111111111010111", 
	 "0111111111010110", 
	 "0111111111010101", 
	 "0111111111010101", 
	 "0111111111010100", 
	 "0111111111010011", 
	 "0111111111010011", 
	 "0111111111010010", 
	 "0111111111010001", 
	 "0111111111010001", 
	 "0111111111010000", 
	 "0111111111001111", 
	 "0111111111001111", 
	 "0111111111001110", 
	 "0111111111001101", 
	 "0111111111001101", 
	 "0111111111001100", 
	 "0111111111001011", 
	 "0111111111001011", 
	 "0111111111001010", 
	 "0111111111001001", 
	 "0111111111001000", 
	 "0111111111001000", 
	 "0111111111000111", 
	 "0111111111000110", 
	 "0111111111000101", 
	 "0111111111000101", 
	 "0111111111000100", 
	 "0111111111000011", 
	 "0111111111000010", 
	 "0111111111000010", 
	 "0111111111000001", 
	 "0111111111000000", 
	 "0111111110111111", 
	 "0111111110111110", 
	 "0111111110111110", 
	 "0111111110111101", 
	 "0111111110111100", 
	 "0111111110111011", 
	 "0111111110111010", 
	 "0111111110111010", 
	 "0111111110111001", 
	 "0111111110111000", 
	 "0111111110110111", 
	 "0111111110110110", 
	 "0111111110110101", 
	 "0111111110110101", 
	 "0111111110110100", 
	 "0111111110110011", 
	 "0111111110110010", 
	 "0111111110110001", 
	 "0111111110110000", 
	 "0111111110101111", 
	 "0111111110101110", 
	 "0111111110101110", 
	 "0111111110101101", 
	 "0111111110101100", 
	 "0111111110101011", 
	 "0111111110101010", 
	 "0111111110101001", 
	 "0111111110101000", 
	 "0111111110100111", 
	 "0111111110100110", 
	 "0111111110100101", 
	 "0111111110100100", 
	 "0111111110100011", 
	 "0111111110100011", 
	 "0111111110100010", 
	 "0111111110100001", 
	 "0111111110100000", 
	 "0111111110011111", 
	 "0111111110011110", 
	 "0111111110011101", 
	 "0111111110011100", 
	 "0111111110011011", 
	 "0111111110011010", 
	 "0111111110011001", 
	 "0111111110011000", 
	 "0111111110010111", 
	 "0111111110010110", 
	 "0111111110010101", 
	 "0111111110010100", 
	 "0111111110010011", 
	 "0111111110010010", 
	 "0111111110010001", 
	 "0111111110010000", 
	 "0111111110001111", 
	 "0111111110001110", 
	 "0111111110001101", 
	 "0111111110001011", 
	 "0111111110001010", 
	 "0111111110001001", 
	 "0111111110001000", 
	 "0111111110000111", 
	 "0111111110000110", 
	 "0111111110000101", 
	 "0111111110000100", 
	 "0111111110000011", 
	 "0111111110000010", 
	 "0111111110000001", 
	 "0111111110000000", 
	 "0111111101111110", 
	 "0111111101111101", 
	 "0111111101111100", 
	 "0111111101111011", 
	 "0111111101111010", 
	 "0111111101111001", 
	 "0111111101111000", 
	 "0111111101110110", 
	 "0111111101110101", 
	 "0111111101110100", 
	 "0111111101110011", 
	 "0111111101110010", 
	 "0111111101110001", 
	 "0111111101101111", 
	 "0111111101101110", 
	 "0111111101101101", 
	 "0111111101101100", 
	 "0111111101101011", 
	 "0111111101101010", 
	 "0111111101101000", 
	 "0111111101100111", 
	 "0111111101100110", 
	 "0111111101100101", 
	 "0111111101100011", 
	 "0111111101100010", 
	 "0111111101100001", 
	 "0111111101100000", 
	 "0111111101011110", 
	 "0111111101011101", 
	 "0111111101011100", 
	 "0111111101011011", 
	 "0111111101011001", 
	 "0111111101011000", 
	 "0111111101010111", 
	 "0111111101010110", 
	 "0111111101010100", 
	 "0111111101010011", 
	 "0111111101010010", 
	 "0111111101010000", 
	 "0111111101001111", 
	 "0111111101001110", 
	 "0111111101001101", 
	 "0111111101001011", 
	 "0111111101001010", 
	 "0111111101001001", 
	 "0111111101000111", 
	 "0111111101000110", 
	 "0111111101000101", 
	 "0111111101000011", 
	 "0111111101000010", 
	 "0111111101000001", 
	 "0111111100111111", 
	 "0111111100111110", 
	 "0111111100111100", 
	 "0111111100111011", 
	 "0111111100111010", 
	 "0111111100111000", 
	 "0111111100110111", 
	 "0111111100110110", 
	 "0111111100110100", 
	 "0111111100110011", 
	 "0111111100110001", 
	 "0111111100110000", 
	 "0111111100101111", 
	 "0111111100101101", 
	 "0111111100101100", 
	 "0111111100101010", 
	 "0111111100101001", 
	 "0111111100100111", 
	 "0111111100100110", 
	 "0111111100100100", 
	 "0111111100100011", 
	 "0111111100100010", 
	 "0111111100100000", 
	 "0111111100011111", 
	 "0111111100011101", 
	 "0111111100011100", 
	 "0111111100011010", 
	 "0111111100011001", 
	 "0111111100010111", 
	 "0111111100010110", 
	 "0111111100010100", 
	 "0111111100010011", 
	 "0111111100010001", 
	 "0111111100010000", 
	 "0111111100001110", 
	 "0111111100001101", 
	 "0111111100001011", 
	 "0111111100001010", 
	 "0111111100001000", 
	 "0111111100000110", 
	 "0111111100000101", 
	 "0111111100000011", 
	 "0111111100000010", 
	 "0111111100000000", 
	 "0111111011111111", 
	 "0111111011111101", 
	 "0111111011111100", 
	 "0111111011111010", 
	 "0111111011111000", 
	 "0111111011110111", 
	 "0111111011110101", 
	 "0111111011110100", 
	 "0111111011110010", 
	 "0111111011110000", 
	 "0111111011101111", 
	 "0111111011101101", 
	 "0111111011101011", 
	 "0111111011101010", 
	 "0111111011101000", 
	 "0111111011100111", 
	 "0111111011100101", 
	 "0111111011100011", 
	 "0111111011100010", 
	 "0111111011100000", 
	 "0111111011011110", 
	 "0111111011011101", 
	 "0111111011011011", 
	 "0111111011011001", 
	 "0111111011011000", 
	 "0111111011010110", 
	 "0111111011010100", 
	 "0111111011010011", 
	 "0111111011010001", 
	 "0111111011001111", 
	 "0111111011001101", 
	 "0111111011001100", 
	 "0111111011001010", 
	 "0111111011001000", 
	 "0111111011000110", 
	 "0111111011000101", 
	 "0111111011000011", 
	 "0111111011000001", 
	 "0111111011000000", 
	 "0111111010111110", 
	 "0111111010111100", 
	 "0111111010111010", 
	 "0111111010111000", 
	 "0111111010110111", 
	 "0111111010110101", 
	 "0111111010110011", 
	 "0111111010110001", 
	 "0111111010110000", 
	 "0111111010101110", 
	 "0111111010101100", 
	 "0111111010101010", 
	 "0111111010101000", 
	 "0111111010100110", 
	 "0111111010100101", 
	 "0111111010100011", 
	 "0111111010100001", 
	 "0111111010011111", 
	 "0111111010011101", 
	 "0111111010011011", 
	 "0111111010011010", 
	 "0111111010011000", 
	 "0111111010010110", 
	 "0111111010010100", 
	 "0111111010010010", 
	 "0111111010010000", 
	 "0111111010001110", 
	 "0111111010001101", 
	 "0111111010001011", 
	 "0111111010001001", 
	 "0111111010000111", 
	 "0111111010000101", 
	 "0111111010000011", 
	 "0111111010000001", 
	 "0111111001111111", 
	 "0111111001111101", 
	 "0111111001111011", 
	 "0111111001111001", 
	 "0111111001111000", 
	 "0111111001110110", 
	 "0111111001110100", 
	 "0111111001110010", 
	 "0111111001110000", 
	 "0111111001101110", 
	 "0111111001101100", 
	 "0111111001101010", 
	 "0111111001101000", 
	 "0111111001100110", 
	 "0111111001100100", 
	 "0111111001100010", 
	 "0111111001100000", 
	 "0111111001011110", 
	 "0111111001011100", 
	 "0111111001011010", 
	 "0111111001011000", 
	 "0111111001010110", 
	 "0111111001010100", 
	 "0111111001010010", 
	 "0111111001010000", 
	 "0111111001001110", 
	 "0111111001001100", 
	 "0111111001001010", 
	 "0111111001001000", 
	 "0111111001000110", 
	 "0111111001000011", 
	 "0111111001000001", 
	 "0111111000111111", 
	 "0111111000111101", 
	 "0111111000111011", 
	 "0111111000111001", 
	 "0111111000110111", 
	 "0111111000110101", 
	 "0111111000110011", 
	 "0111111000110001", 
	 "0111111000101111", 
	 "0111111000101101", 
	 "0111111000101010", 
	 "0111111000101000", 
	 "0111111000100110", 
	 "0111111000100100", 
	 "0111111000100010", 
	 "0111111000100000", 
	 "0111111000011110", 
	 "0111111000011011", 
	 "0111111000011001", 
	 "0111111000010111", 
	 "0111111000010101", 
	 "0111111000010011", 
	 "0111111000010001", 
	 "0111111000001110", 
	 "0111111000001100", 
	 "0111111000001010", 
	 "0111111000001000", 
	 "0111111000000110", 
	 "0111111000000011", 
	 "0111111000000001", 
	 "0111110111111111", 
	 "0111110111111101", 
	 "0111110111111011", 
	 "0111110111111000", 
	 "0111110111110110", 
	 "0111110111110100", 
	 "0111110111110010", 
	 "0111110111101111", 
	 "0111110111101101", 
	 "0111110111101011", 
	 "0111110111101001", 
	 "0111110111100110", 
	 "0111110111100100", 
	 "0111110111100010", 
	 "0111110111100000", 
	 "0111110111011101", 
	 "0111110111011011", 
	 "0111110111011001", 
	 "0111110111010110", 
	 "0111110111010100", 
	 "0111110111010010", 
	 "0111110111001111", 
	 "0111110111001101", 
	 "0111110111001011", 
	 "0111110111001001", 
	 "0111110111000110", 
	 "0111110111000100", 
	 "0111110111000010", 
	 "0111110110111111", 
	 "0111110110111101", 
	 "0111110110111010", 
	 "0111110110111000", 
	 "0111110110110110", 
	 "0111110110110011", 
	 "0111110110110001", 
	 "0111110110101111", 
	 "0111110110101100", 
	 "0111110110101010", 
	 "0111110110100111", 
	 "0111110110100101", 
	 "0111110110100011", 
	 "0111110110100000", 
	 "0111110110011110", 
	 "0111110110011011", 
	 "0111110110011001", 
	 "0111110110010111", 
	 "0111110110010100", 
	 "0111110110010010", 
	 "0111110110001111", 
	 "0111110110001101", 
	 "0111110110001010", 
	 "0111110110001000", 
	 "0111110110000101", 
	 "0111110110000011", 
	 "0111110110000001", 
	 "0111110101111110", 
	 "0111110101111100", 
	 "0111110101111001", 
	 "0111110101110111", 
	 "0111110101110100", 
	 "0111110101110010", 
	 "0111110101101111", 
	 "0111110101101101", 
	 "0111110101101010", 
	 "0111110101101000", 
	 "0111110101100101", 
	 "0111110101100011", 
	 "0111110101100000", 
	 "0111110101011101", 
	 "0111110101011011", 
	 "0111110101011000", 
	 "0111110101010110", 
	 "0111110101010011", 
	 "0111110101010001", 
	 "0111110101001110", 
	 "0111110101001100", 
	 "0111110101001001", 
	 "0111110101000110", 
	 "0111110101000100", 
	 "0111110101000001", 
	 "0111110100111111", 
	 "0111110100111100", 
	 "0111110100111010", 
	 "0111110100110111", 
	 "0111110100110100", 
	 "0111110100110010", 
	 "0111110100101111", 
	 "0111110100101100", 
	 "0111110100101010", 
	 "0111110100100111", 
	 "0111110100100101", 
	 "0111110100100010", 
	 "0111110100011111", 
	 "0111110100011101", 
	 "0111110100011010", 
	 "0111110100010111", 
	 "0111110100010101", 
	 "0111110100010010", 
	 "0111110100001111", 
	 "0111110100001101", 
	 "0111110100001010", 
	 "0111110100000111", 
	 "0111110100000101", 
	 "0111110100000010", 
	 "0111110011111111", 
	 "0111110011111100", 
	 "0111110011111010", 
	 "0111110011110111", 
	 "0111110011110100", 
	 "0111110011110010", 
	 "0111110011101111", 
	 "0111110011101100", 
	 "0111110011101001", 
	 "0111110011100111", 
	 "0111110011100100", 
	 "0111110011100001", 
	 "0111110011011110", 
	 "0111110011011100", 
	 "0111110011011001", 
	 "0111110011010110", 
	 "0111110011010011", 
	 "0111110011010000", 
	 "0111110011001110", 
	 "0111110011001011", 
	 "0111110011001000", 
	 "0111110011000101", 
	 "0111110011000010", 
	 "0111110011000000", 
	 "0111110010111101", 
	 "0111110010111010", 
	 "0111110010110111", 
	 "0111110010110100", 
	 "0111110010110001", 
	 "0111110010101111", 
	 "0111110010101100", 
	 "0111110010101001", 
	 "0111110010100110", 
	 "0111110010100011", 
	 "0111110010100000", 
	 "0111110010011110", 
	 "0111110010011011", 
	 "0111110010011000", 
	 "0111110010010101", 
	 "0111110010010010", 
	 "0111110010001111", 
	 "0111110010001100", 
	 "0111110010001001", 
	 "0111110010000110", 
	 "0111110010000011", 
	 "0111110010000001", 
	 "0111110001111110", 
	 "0111110001111011", 
	 "0111110001111000", 
	 "0111110001110101", 
	 "0111110001110010", 
	 "0111110001101111", 
	 "0111110001101100", 
	 "0111110001101001", 
	 "0111110001100110", 
	 "0111110001100011", 
	 "0111110001100000", 
	 "0111110001011101", 
	 "0111110001011010", 
	 "0111110001010111", 
	 "0111110001010100", 
	 "0111110001010001", 
	 "0111110001001110", 
	 "0111110001001011", 
	 "0111110001001000", 
	 "0111110001000101", 
	 "0111110001000010", 
	 "0111110000111111", 
	 "0111110000111100", 
	 "0111110000111001", 
	 "0111110000110110", 
	 "0111110000110011", 
	 "0111110000110000", 
	 "0111110000101101", 
	 "0111110000101010", 
	 "0111110000100111", 
	 "0111110000100100", 
	 "0111110000100001", 
	 "0111110000011110", 
	 "0111110000011011", 
	 "0111110000011000", 
	 "0111110000010100", 
	 "0111110000010001", 
	 "0111110000001110", 
	 "0111110000001011", 
	 "0111110000001000", 
	 "0111110000000101", 
	 "0111110000000010", 
	 "0111101111111111", 
	 "0111101111111100", 
	 "0111101111111001", 
	 "0111101111110101", 
	 "0111101111110010", 
	 "0111101111101111", 
	 "0111101111101100", 
	 "0111101111101001", 
	 "0111101111100110", 
	 "0111101111100011", 
	 "0111101111011111", 
	 "0111101111011100", 
	 "0111101111011001", 
	 "0111101111010110", 
	 "0111101111010011", 
	 "0111101111001111", 
	 "0111101111001100", 
	 "0111101111001001", 
	 "0111101111000110", 
	 "0111101111000011", 
	 "0111101110111111", 
	 "0111101110111100", 
	 "0111101110111001", 
	 "0111101110110110", 
	 "0111101110110011", 
	 "0111101110101111", 
	 "0111101110101100", 
	 "0111101110101001", 
	 "0111101110100110", 
	 "0111101110100010", 
	 "0111101110011111", 
	 "0111101110011100", 
	 "0111101110011001", 
	 "0111101110010101", 
	 "0111101110010010", 
	 "0111101110001111", 
	 "0111101110001011", 
	 "0111101110001000", 
	 "0111101110000101", 
	 "0111101110000010", 
	 "0111101101111110", 
	 "0111101101111011", 
	 "0111101101111000", 
	 "0111101101110100", 
	 "0111101101110001", 
	 "0111101101101110", 
	 "0111101101101010", 
	 "0111101101100111", 
	 "0111101101100100", 
	 "0111101101100000", 
	 "0111101101011101", 
	 "0111101101011010", 
	 "0111101101010110", 
	 "0111101101010011", 
	 "0111101101010000", 
	 "0111101101001100", 
	 "0111101101001001", 
	 "0111101101000101", 
	 "0111101101000010", 
	 "0111101100111111", 
	 "0111101100111011", 
	 "0111101100111000", 
	 "0111101100110100", 
	 "0111101100110001", 
	 "0111101100101110", 
	 "0111101100101010", 
	 "0111101100100111", 
	 "0111101100100011", 
	 "0111101100100000", 
	 "0111101100011100", 
	 "0111101100011001", 
	 "0111101100010110", 
	 "0111101100010010", 
	 "0111101100001111", 
	 "0111101100001011", 
	 "0111101100001000", 
	 "0111101100000100", 
	 "0111101100000001", 
	 "0111101011111101", 
	 "0111101011111010", 
	 "0111101011110110", 
	 "0111101011110011", 
	 "0111101011101111", 
	 "0111101011101100", 
	 "0111101011101000", 
	 "0111101011100101", 
	 "0111101011100001", 
	 "0111101011011110", 
	 "0111101011011010", 
	 "0111101011010111", 
	 "0111101011010011", 
	 "0111101011010000", 
	 "0111101011001100", 
	 "0111101011001001", 
	 "0111101011000101", 
	 "0111101011000001", 
	 "0111101010111110", 
	 "0111101010111010", 
	 "0111101010110111", 
	 "0111101010110011", 
	 "0111101010110000", 
	 "0111101010101100", 
	 "0111101010101000", 
	 "0111101010100101", 
	 "0111101010100001", 
	 "0111101010011110", 
	 "0111101010011010", 
	 "0111101010010110", 
	 "0111101010010011", 
	 "0111101010001111", 
	 "0111101010001100", 
	 "0111101010001000", 
	 "0111101010000100", 
	 "0111101010000001", 
	 "0111101001111101", 
	 "0111101001111001", 
	 "0111101001110110", 
	 "0111101001110010", 
	 "0111101001101110", 
	 "0111101001101011", 
	 "0111101001100111", 
	 "0111101001100011", 
	 "0111101001100000", 
	 "0111101001011100", 
	 "0111101001011000", 
	 "0111101001010101", 
	 "0111101001010001", 
	 "0111101001001101", 
	 "0111101001001001", 
	 "0111101001000110", 
	 "0111101001000010", 
	 "0111101000111110", 
	 "0111101000111011", 
	 "0111101000110111", 
	 "0111101000110011", 
	 "0111101000101111", 
	 "0111101000101100", 
	 "0111101000101000", 
	 "0111101000100100", 
	 "0111101000100000", 
	 "0111101000011101", 
	 "0111101000011001", 
	 "0111101000010101", 
	 "0111101000010001", 
	 "0111101000001110", 
	 "0111101000001010", 
	 "0111101000000110", 
	 "0111101000000010", 
	 "0111100111111110", 
	 "0111100111111011", 
	 "0111100111110111", 
	 "0111100111110011", 
	 "0111100111101111", 
	 "0111100111101011", 
	 "0111100111100111", 
	 "0111100111100100", 
	 "0111100111100000", 
	 "0111100111011100", 
	 "0111100111011000", 
	 "0111100111010100", 
	 "0111100111010000", 
	 "0111100111001100", 
	 "0111100111001001", 
	 "0111100111000101", 
	 "0111100111000001", 
	 "0111100110111101", 
	 "0111100110111001", 
	 "0111100110110101", 
	 "0111100110110001", 
	 "0111100110101101", 
	 "0111100110101010", 
	 "0111100110100110", 
	 "0111100110100010", 
	 "0111100110011110", 
	 "0111100110011010", 
	 "0111100110010110", 
	 "0111100110010010", 
	 "0111100110001110", 
	 "0111100110001010", 
	 "0111100110000110", 
	 "0111100110000010", 
	 "0111100101111110", 
	 "0111100101111010", 
	 "0111100101110110", 
	 "0111100101110010", 
	 "0111100101101110", 
	 "0111100101101010", 
	 "0111100101100110", 
	 "0111100101100010", 
	 "0111100101011111", 
	 "0111100101011011", 
	 "0111100101010111", 
	 "0111100101010011", 
	 "0111100101001110", 
	 "0111100101001010", 
	 "0111100101000110", 
	 "0111100101000010", 
	 "0111100100111110", 
	 "0111100100111010", 
	 "0111100100110110", 
	 "0111100100110010", 
	 "0111100100101110", 
	 "0111100100101010", 
	 "0111100100100110", 
	 "0111100100100010", 
	 "0111100100011110", 
	 "0111100100011010", 
	 "0111100100010110", 
	 "0111100100010010", 
	 "0111100100001110", 
	 "0111100100001010", 
	 "0111100100000110", 
	 "0111100100000001", 
	 "0111100011111101", 
	 "0111100011111001", 
	 "0111100011110101", 
	 "0111100011110001", 
	 "0111100011101101", 
	 "0111100011101001", 
	 "0111100011100101", 
	 "0111100011100001", 
	 "0111100011011100", 
	 "0111100011011000", 
	 "0111100011010100", 
	 "0111100011010000", 
	 "0111100011001100", 
	 "0111100011001000", 
	 "0111100011000100", 
	 "0111100010111111", 
	 "0111100010111011", 
	 "0111100010110111", 
	 "0111100010110011", 
	 "0111100010101111", 
	 "0111100010101010", 
	 "0111100010100110", 
	 "0111100010100010", 
	 "0111100010011110", 
	 "0111100010011010", 
	 "0111100010010101", 
	 "0111100010010001", 
	 "0111100010001101", 
	 "0111100010001001", 
	 "0111100010000101", 
	 "0111100010000000", 
	 "0111100001111100", 
	 "0111100001111000", 
	 "0111100001110100", 
	 "0111100001101111", 
	 "0111100001101011", 
	 "0111100001100111", 
	 "0111100001100011", 
	 "0111100001011110", 
	 "0111100001011010", 
	 "0111100001010110", 
	 "0111100001010001", 
	 "0111100001001101", 
	 "0111100001001001", 
	 "0111100001000101", 
	 "0111100001000000", 
	 "0111100000111100", 
	 "0111100000111000", 
	 "0111100000110011", 
	 "0111100000101111", 
	 "0111100000101011", 
	 "0111100000100110", 
	 "0111100000100010", 
	 "0111100000011110", 
	 "0111100000011001", 
	 "0111100000010101", 
	 "0111100000010001", 
	 "0111100000001100", 
	 "0111100000001000", 
	 "0111100000000011", 
	 "0111011111111111", 
	 "0111011111111011", 
	 "0111011111110110", 
	 "0111011111110010", 
	 "0111011111101110", 
	 "0111011111101001", 
	 "0111011111100101", 
	 "0111011111100000", 
	 "0111011111011100", 
	 "0111011111011000", 
	 "0111011111010011", 
	 "0111011111001111", 
	 "0111011111001010", 
	 "0111011111000110", 
	 "0111011111000001", 
	 "0111011110111101", 
	 "0111011110111001", 
	 "0111011110110100", 
	 "0111011110110000", 
	 "0111011110101011", 
	 "0111011110100111", 
	 "0111011110100010", 
	 "0111011110011110", 
	 "0111011110011001", 
	 "0111011110010101", 
	 "0111011110010000", 
	 "0111011110001100", 
	 "0111011110000111", 
	 "0111011110000011", 
	 "0111011101111110", 
	 "0111011101111010", 
	 "0111011101110101", 
	 "0111011101110001", 
	 "0111011101101100", 
	 "0111011101101000", 
	 "0111011101100011", 
	 "0111011101011111", 
	 "0111011101011010", 
	 "0111011101010110", 
	 "0111011101010001", 
	 "0111011101001101", 
	 "0111011101001000", 
	 "0111011101000011", 
	 "0111011100111111", 
	 "0111011100111010", 
	 "0111011100110110", 
	 "0111011100110001", 
	 "0111011100101101", 
	 "0111011100101000", 
	 "0111011100100011", 
	 "0111011100011111", 
	 "0111011100011010", 
	 "0111011100010110", 
	 "0111011100010001", 
	 "0111011100001100", 
	 "0111011100001000", 
	 "0111011100000011", 
	 "0111011011111110", 
	 "0111011011111010", 
	 "0111011011110101", 
	 "0111011011110001", 
	 "0111011011101100", 
	 "0111011011100111", 
	 "0111011011100011", 
	 "0111011011011110", 
	 "0111011011011001", 
	 "0111011011010101", 
	 "0111011011010000", 
	 "0111011011001011", 
	 "0111011011000111", 
	 "0111011011000010", 
	 "0111011010111101", 
	 "0111011010111001", 
	 "0111011010110100", 
	 "0111011010101111", 
	 "0111011010101010", 
	 "0111011010100110", 
	 "0111011010100001", 
	 "0111011010011100", 
	 "0111011010011000", 
	 "0111011010010011", 
	 "0111011010001110", 
	 "0111011010001001", 
	 "0111011010000101", 
	 "0111011010000000", 
	 "0111011001111011", 
	 "0111011001110110", 
	 "0111011001110010", 
	 "0111011001101101", 
	 "0111011001101000", 
	 "0111011001100011", 
	 "0111011001011110", 
	 "0111011001011010", 
	 "0111011001010101", 
	 "0111011001010000", 
	 "0111011001001011", 
	 "0111011001000110", 
	 "0111011001000010", 
	 "0111011000111101", 
	 "0111011000111000", 
	 "0111011000110011", 
	 "0111011000101110", 
	 "0111011000101010", 
	 "0111011000100101", 
	 "0111011000100000", 
	 "0111011000011011", 
	 "0111011000010110", 
	 "0111011000010001", 
	 "0111011000001101", 
	 "0111011000001000", 
	 "0111011000000011", 
	 "0111010111111110", 
	 "0111010111111001", 
	 "0111010111110100", 
	 "0111010111101111", 
	 "0111010111101010", 
	 "0111010111100110", 
	 "0111010111100001", 
	 "0111010111011100", 
	 "0111010111010111", 
	 "0111010111010010", 
	 "0111010111001101", 
	 "0111010111001000", 
	 "0111010111000011", 
	 "0111010110111110", 
	 "0111010110111001", 
	 "0111010110110100", 
	 "0111010110101111", 
	 "0111010110101010", 
	 "0111010110100110", 
	 "0111010110100001", 
	 "0111010110011100", 
	 "0111010110010111", 
	 "0111010110010010", 
	 "0111010110001101", 
	 "0111010110001000", 
	 "0111010110000011", 
	 "0111010101111110", 
	 "0111010101111001", 
	 "0111010101110100", 
	 "0111010101101111", 
	 "0111010101101010", 
	 "0111010101100101", 
	 "0111010101100000", 
	 "0111010101011011", 
	 "0111010101010110", 
	 "0111010101010001", 
	 "0111010101001100", 
	 "0111010101000111", 
	 "0111010101000010", 
	 "0111010100111101", 
	 "0111010100111000", 
	 "0111010100110010", 
	 "0111010100101101", 
	 "0111010100101000", 
	 "0111010100100011", 
	 "0111010100011110", 
	 "0111010100011001", 
	 "0111010100010100", 
	 "0111010100001111", 
	 "0111010100001010", 
	 "0111010100000101", 
	 "0111010100000000", 
	 "0111010011111011", 
	 "0111010011110110", 
	 "0111010011110000", 
	 "0111010011101011", 
	 "0111010011100110", 
	 "0111010011100001", 
	 "0111010011011100", 
	 "0111010011010111", 
	 "0111010011010010", 
	 "0111010011001101", 
	 "0111010011000111", 
	 "0111010011000010", 
	 "0111010010111101", 
	 "0111010010111000", 
	 "0111010010110011", 
	 "0111010010101110", 
	 "0111010010101000", 
	 "0111010010100011", 
	 "0111010010011110", 
	 "0111010010011001", 
	 "0111010010010100", 
	 "0111010010001111", 
	 "0111010010001001", 
	 "0111010010000100", 
	 "0111010001111111", 
	 "0111010001111010", 
	 "0111010001110101", 
	 "0111010001101111", 
	 "0111010001101010", 
	 "0111010001100101", 
	 "0111010001100000", 
	 "0111010001011010", 
	 "0111010001010101", 
	 "0111010001010000", 
	 "0111010001001011", 
	 "0111010001000101", 
	 "0111010001000000", 
	 "0111010000111011", 
	 "0111010000110110", 
	 "0111010000110000", 
	 "0111010000101011", 
	 "0111010000100110", 
	 "0111010000100001", 
	 "0111010000011011", 
	 "0111010000010110", 
	 "0111010000010001", 
	 "0111010000001011", 
	 "0111010000000110", 
	 "0111010000000001", 
	 "0111001111111011", 
	 "0111001111110110", 
	 "0111001111110001", 
	 "0111001111101011", 
	 "0111001111100110", 
	 "0111001111100001", 
	 "0111001111011011", 
	 "0111001111010110", 
	 "0111001111010001", 
	 "0111001111001011", 
	 "0111001111000110", 
	 "0111001111000001", 
	 "0111001110111011", 
	 "0111001110110110", 
	 "0111001110110001", 
	 "0111001110101011", 
	 "0111001110100110", 
	 "0111001110100000", 
	 "0111001110011011", 
	 "0111001110010110", 
	 "0111001110010000", 
	 "0111001110001011", 
	 "0111001110000101", 
	 "0111001110000000", 
	 "0111001101111011", 
	 "0111001101110101", 
	 "0111001101110000", 
	 "0111001101101010", 
	 "0111001101100101", 
	 "0111001101011111", 
	 "0111001101011010", 
	 "0111001101010101", 
	 "0111001101001111", 
	 "0111001101001010", 
	 "0111001101000100", 
	 "0111001100111111", 
	 "0111001100111001", 
	 "0111001100110100", 
	 "0111001100101110", 
	 "0111001100101001", 
	 "0111001100100011", 
	 "0111001100011110", 
	 "0111001100011000", 
	 "0111001100010011", 
	 "0111001100001101", 
	 "0111001100001000", 
	 "0111001100000010", 
	 "0111001011111101", 
	 "0111001011110111", 
	 "0111001011110010", 
	 "0111001011101100", 
	 "0111001011100111", 
	 "0111001011100001", 
	 "0111001011011100", 
	 "0111001011010110", 
	 "0111001011010000", 
	 "0111001011001011", 
	 "0111001011000101", 
	 "0111001011000000", 
	 "0111001010111010", 
	 "0111001010110101", 
	 "0111001010101111", 
	 "0111001010101001", 
	 "0111001010100100", 
	 "0111001010011110", 
	 "0111001010011001", 
	 "0111001010010011", 
	 "0111001010001101", 
	 "0111001010001000", 
	 "0111001010000010", 
	 "0111001001111101", 
	 "0111001001110111", 
	 "0111001001110001", 
	 "0111001001101100", 
	 "0111001001100110", 
	 "0111001001100000", 
	 "0111001001011011", 
	 "0111001001010101", 
	 "0111001001010000", 
	 "0111001001001010", 
	 "0111001001000100", 
	 "0111001000111111", 
	 "0111001000111001", 
	 "0111001000110011", 
	 "0111001000101110", 
	 "0111001000101000", 
	 "0111001000100010", 
	 "0111001000011100", 
	 "0111001000010111", 
	 "0111001000010001", 
	 "0111001000001011", 
	 "0111001000000110", 
	 "0111001000000000", 
	 "0111000111111010", 
	 "0111000111110101", 
	 "0111000111101111", 
	 "0111000111101001", 
	 "0111000111100011", 
	 "0111000111011110", 
	 "0111000111011000", 
	 "0111000111010010", 
	 "0111000111001100", 
	 "0111000111000111", 
	 "0111000111000001", 
	 "0111000110111011", 
	 "0111000110110101", 
	 "0111000110110000", 
	 "0111000110101010", 
	 "0111000110100100", 
	 "0111000110011110", 
	 "0111000110011000", 
	 "0111000110010011", 
	 "0111000110001101", 
	 "0111000110000111", 
	 "0111000110000001", 
	 "0111000101111011", 
	 "0111000101110110", 
	 "0111000101110000", 
	 "0111000101101010", 
	 "0111000101100100", 
	 "0111000101011110", 
	 "0111000101011000", 
	 "0111000101010011", 
	 "0111000101001101", 
	 "0111000101000111", 
	 "0111000101000001", 
	 "0111000100111011", 
	 "0111000100110101", 
	 "0111000100101111", 
	 "0111000100101010", 
	 "0111000100100100", 
	 "0111000100011110", 
	 "0111000100011000", 
	 "0111000100010010", 
	 "0111000100001100", 
	 "0111000100000110", 
	 "0111000100000000", 
	 "0111000011111010", 
	 "0111000011110101", 
	 "0111000011101111", 
	 "0111000011101001", 
	 "0111000011100011", 
	 "0111000011011101", 
	 "0111000011010111", 
	 "0111000011010001", 
	 "0111000011001011", 
	 "0111000011000101", 
	 "0111000010111111", 
	 "0111000010111001", 
	 "0111000010110011", 
	 "0111000010101101", 
	 "0111000010100111", 
	 "0111000010100001", 
	 "0111000010011011", 
	 "0111000010010101", 
	 "0111000010001111", 
	 "0111000010001001", 
	 "0111000010000011", 
	 "0111000001111101", 
	 "0111000001110111", 
	 "0111000001110001", 
	 "0111000001101011", 
	 "0111000001100101", 
	 "0111000001011111", 
	 "0111000001011001", 
	 "0111000001010011", 
	 "0111000001001101", 
	 "0111000001000111", 
	 "0111000001000001", 
	 "0111000000111011", 
	 "0111000000110101", 
	 "0111000000101111", 
	 "0111000000101001", 
	 "0111000000100011", 
	 "0111000000011101", 
	 "0111000000010111", 
	 "0111000000010001", 
	 "0111000000001011", 
	 "0111000000000101", 
	 "0110111111111111", 
	 "0110111111111001", 
	 "0110111111110010", 
	 "0110111111101100", 
	 "0110111111100110", 
	 "0110111111100000", 
	 "0110111111011010", 
	 "0110111111010100", 
	 "0110111111001110", 
	 "0110111111001000", 
	 "0110111111000010", 
	 "0110111110111011", 
	 "0110111110110101", 
	 "0110111110101111", 
	 "0110111110101001", 
	 "0110111110100011", 
	 "0110111110011101", 
	 "0110111110010111", 
	 "0110111110010000", 
	 "0110111110001010", 
	 "0110111110000100", 
	 "0110111101111110", 
	 "0110111101111000", 
	 "0110111101110010", 
	 "0110111101101011", 
	 "0110111101100101", 
	 "0110111101011111", 
	 "0110111101011001", 
	 "0110111101010011", 
	 "0110111101001100", 
	 "0110111101000110", 
	 "0110111101000000", 
	 "0110111100111010", 
	 "0110111100110100", 
	 "0110111100101101", 
	 "0110111100100111", 
	 "0110111100100001", 
	 "0110111100011011", 
	 "0110111100010100", 
	 "0110111100001110", 
	 "0110111100001000", 
	 "0110111100000010", 
	 "0110111011111011", 
	 "0110111011110101", 
	 "0110111011101111", 
	 "0110111011101001", 
	 "0110111011100010", 
	 "0110111011011100", 
	 "0110111011010110", 
	 "0110111011001111", 
	 "0110111011001001", 
	 "0110111011000011", 
	 "0110111010111101", 
	 "0110111010110110", 
	 "0110111010110000", 
	 "0110111010101010", 
	 "0110111010100011", 
	 "0110111010011101", 
	 "0110111010010111", 
	 "0110111010010000", 
	 "0110111010001010", 
	 "0110111010000100", 
	 "0110111001111101", 
	 "0110111001110111", 
	 "0110111001110001", 
	 "0110111001101010", 
	 "0110111001100100", 
	 "0110111001011110", 
	 "0110111001010111", 
	 "0110111001010001", 
	 "0110111001001010", 
	 "0110111001000100", 
	 "0110111000111110", 
	 "0110111000110111", 
	 "0110111000110001", 
	 "0110111000101010", 
	 "0110111000100100", 
	 "0110111000011110", 
	 "0110111000010111", 
	 "0110111000010001", 
	 "0110111000001010", 
	 "0110111000000100", 
	 "0110110111111110", 
	 "0110110111110111", 
	 "0110110111110001", 
	 "0110110111101010", 
	 "0110110111100100", 
	 "0110110111011101", 
	 "0110110111010111", 
	 "0110110111010001", 
	 "0110110111001010", 
	 "0110110111000100", 
	 "0110110110111101", 
	 "0110110110110111", 
	 "0110110110110000", 
	 "0110110110101010", 
	 "0110110110100011", 
	 "0110110110011101", 
	 "0110110110010110", 
	 "0110110110010000", 
	 "0110110110001001", 
	 "0110110110000011", 
	 "0110110101111100", 
	 "0110110101110110", 
	 "0110110101101111", 
	 "0110110101101001", 
	 "0110110101100010", 
	 "0110110101011100", 
	 "0110110101010101", 
	 "0110110101001111", 
	 "0110110101001000", 
	 "0110110101000001", 
	 "0110110100111011", 
	 "0110110100110100", 
	 "0110110100101110", 
	 "0110110100100111", 
	 "0110110100100001", 
	 "0110110100011010", 
	 "0110110100010100", 
	 "0110110100001101", 
	 "0110110100000110", 
	 "0110110100000000", 
	 "0110110011111001", 
	 "0110110011110011", 
	 "0110110011101100", 
	 "0110110011100101", 
	 "0110110011011111", 
	 "0110110011011000", 
	 "0110110011010010", 
	 "0110110011001011", 
	 "0110110011000100", 
	 "0110110010111110", 
	 "0110110010110111", 
	 "0110110010110000", 
	 "0110110010101010", 
	 "0110110010100011", 
	 "0110110010011101", 
	 "0110110010010110", 
	 "0110110010001111", 
	 "0110110010001001", 
	 "0110110010000010", 
	 "0110110001111011", 
	 "0110110001110101", 
	 "0110110001101110", 
	 "0110110001100111", 
	 "0110110001100001", 
	 "0110110001011010", 
	 "0110110001010011", 
	 "0110110001001100", 
	 "0110110001000110", 
	 "0110110000111111", 
	 "0110110000111000", 
	 "0110110000110010", 
	 "0110110000101011", 
	 "0110110000100100", 
	 "0110110000011101", 
	 "0110110000010111", 
	 "0110110000010000", 
	 "0110110000001001", 
	 "0110110000000010", 
	 "0110101111111100", 
	 "0110101111110101", 
	 "0110101111101110", 
	 "0110101111100111", 
	 "0110101111100001", 
	 "0110101111011010", 
	 "0110101111010011", 
	 "0110101111001100", 
	 "0110101111000110", 
	 "0110101110111111", 
	 "0110101110111000", 
	 "0110101110110001", 
	 "0110101110101010", 
	 "0110101110100100", 
	 "0110101110011101", 
	 "0110101110010110", 
	 "0110101110001111", 
	 "0110101110001000", 
	 "0110101110000010", 
	 "0110101101111011", 
	 "0110101101110100", 
	 "0110101101101101", 
	 "0110101101100110", 
	 "0110101101011111", 
	 "0110101101011001", 
	 "0110101101010010", 
	 "0110101101001011", 
	 "0110101101000100", 
	 "0110101100111101", 
	 "0110101100110110", 
	 "0110101100110000", 
	 "0110101100101001", 
	 "0110101100100010", 
	 "0110101100011011", 
	 "0110101100010100", 
	 "0110101100001101", 
	 "0110101100000110", 
	 "0110101011111111", 
	 "0110101011111000", 
	 "0110101011110010", 
	 "0110101011101011", 
	 "0110101011100100", 
	 "0110101011011101", 
	 "0110101011010110", 
	 "0110101011001111", 
	 "0110101011001000", 
	 "0110101011000001", 
	 "0110101010111010", 
	 "0110101010110011", 
	 "0110101010101100", 
	 "0110101010100101", 
	 "0110101010011110", 
	 "0110101010010111", 
	 "0110101010010000", 
	 "0110101010001001", 
	 "0110101010000011", 
	 "0110101001111100", 
	 "0110101001110101", 
	 "0110101001101110", 
	 "0110101001100111", 
	 "0110101001100000", 
	 "0110101001011001", 
	 "0110101001010010", 
	 "0110101001001011", 
	 "0110101001000100", 
	 "0110101000111101", 
	 "0110101000110110", 
	 "0110101000101111", 
	 "0110101000101000", 
	 "0110101000100001", 
	 "0110101000011010", 
	 "0110101000010010", 
	 "0110101000001011", 
	 "0110101000000100", 
	 "0110100111111101", 
	 "0110100111110110", 
	 "0110100111101111", 
	 "0110100111101000", 
	 "0110100111100001", 
	 "0110100111011010", 
	 "0110100111010011", 
	 "0110100111001100", 
	 "0110100111000101", 
	 "0110100110111110", 
	 "0110100110110111", 
	 "0110100110110000", 
	 "0110100110101001", 
	 "0110100110100001", 
	 "0110100110011010", 
	 "0110100110010011", 
	 "0110100110001100", 
	 "0110100110000101", 
	 "0110100101111110", 
	 "0110100101110111", 
	 "0110100101110000", 
	 "0110100101101001", 
	 "0110100101100001", 
	 "0110100101011010", 
	 "0110100101010011", 
	 "0110100101001100", 
	 "0110100101000101", 
	 "0110100100111110", 
	 "0110100100110111", 
	 "0110100100101111", 
	 "0110100100101000", 
	 "0110100100100001", 
	 "0110100100011010", 
	 "0110100100010011", 
	 "0110100100001100", 
	 "0110100100000100", 
	 "0110100011111101", 
	 "0110100011110110", 
	 "0110100011101111", 
	 "0110100011101000", 
	 "0110100011100000", 
	 "0110100011011001", 
	 "0110100011010010", 
	 "0110100011001011", 
	 "0110100011000100", 
	 "0110100010111100", 
	 "0110100010110101", 
	 "0110100010101110", 
	 "0110100010100111", 
	 "0110100010011111", 
	 "0110100010011000", 
	 "0110100010010001", 
	 "0110100010001010", 
	 "0110100010000010", 
	 "0110100001111011", 
	 "0110100001110100", 
	 "0110100001101101", 
	 "0110100001100101", 
	 "0110100001011110", 
	 "0110100001010111", 
	 "0110100001010000", 
	 "0110100001001000", 
	 "0110100001000001", 
	 "0110100000111010", 
	 "0110100000110010", 
	 "0110100000101011", 
	 "0110100000100100", 
	 "0110100000011100", 
	 "0110100000010101", 
	 "0110100000001110", 
	 "0110100000000110", 
	 "0110011111111111", 
	 "0110011111111000", 
	 "0110011111110000", 
	 "0110011111101001", 
	 "0110011111100010", 
	 "0110011111011010", 
	 "0110011111010011", 
	 "0110011111001100", 
	 "0110011111000100", 
	 "0110011110111101", 
	 "0110011110110110", 
	 "0110011110101110", 
	 "0110011110100111", 
	 "0110011110100000", 
	 "0110011110011000", 
	 "0110011110010001", 
	 "0110011110001001", 
	 "0110011110000010", 
	 "0110011101111011", 
	 "0110011101110011", 
	 "0110011101101100", 
	 "0110011101100100", 
	 "0110011101011101", 
	 "0110011101010110", 
	 "0110011101001110", 
	 "0110011101000111", 
	 "0110011100111111", 
	 "0110011100111000", 
	 "0110011100110000", 
	 "0110011100101001", 
	 "0110011100100010", 
	 "0110011100011010", 
	 "0110011100010011", 
	 "0110011100001011", 
	 "0110011100000100", 
	 "0110011011111100", 
	 "0110011011110101", 
	 "0110011011101101", 
	 "0110011011100110", 
	 "0110011011011110", 
	 "0110011011010111", 
	 "0110011011010000", 
	 "0110011011001000", 
	 "0110011011000001", 
	 "0110011010111001", 
	 "0110011010110010", 
	 "0110011010101010", 
	 "0110011010100011", 
	 "0110011010011011", 
	 "0110011010010011", 
	 "0110011010001100", 
	 "0110011010000100", 
	 "0110011001111101", 
	 "0110011001110101", 
	 "0110011001101110", 
	 "0110011001100110", 
	 "0110011001011111", 
	 "0110011001010111", 
	 "0110011001010000", 
	 "0110011001001000", 
	 "0110011001000001", 
	 "0110011000111001", 
	 "0110011000110001", 
	 "0110011000101010", 
	 "0110011000100010", 
	 "0110011000011011", 
	 "0110011000010011", 
	 "0110011000001100", 
	 "0110011000000100", 
	 "0110010111111100", 
	 "0110010111110101", 
	 "0110010111101101", 
	 "0110010111100110", 
	 "0110010111011110", 
	 "0110010111010110", 
	 "0110010111001111", 
	 "0110010111000111", 
	 "0110010111000000", 
	 "0110010110111000", 
	 "0110010110110000", 
	 "0110010110101001", 
	 "0110010110100001", 
	 "0110010110011001", 
	 "0110010110010010", 
	 "0110010110001010", 
	 "0110010110000010", 
	 "0110010101111011", 
	 "0110010101110011", 
	 "0110010101101011", 
	 "0110010101100100", 
	 "0110010101011100", 
	 "0110010101010100", 
	 "0110010101001101", 
	 "0110010101000101", 
	 "0110010100111101", 
	 "0110010100110110", 
	 "0110010100101110", 
	 "0110010100100110", 
	 "0110010100011111", 
	 "0110010100010111", 
	 "0110010100001111", 
	 "0110010100000111", 
	 "0110010100000000", 
	 "0110010011111000", 
	 "0110010011110000", 
	 "0110010011101001", 
	 "0110010011100001", 
	 "0110010011011001", 
	 "0110010011010001", 
	 "0110010011001010", 
	 "0110010011000010", 
	 "0110010010111010", 
	 "0110010010110010", 
	 "0110010010101011", 
	 "0110010010100011", 
	 "0110010010011011", 
	 "0110010010010011", 
	 "0110010010001011", 
	 "0110010010000100", 
	 "0110010001111100", 
	 "0110010001110100", 
	 "0110010001101100", 
	 "0110010001100101", 
	 "0110010001011101", 
	 "0110010001010101", 
	 "0110010001001101", 
	 "0110010001000101", 
	 "0110010000111110", 
	 "0110010000110110", 
	 "0110010000101110", 
	 "0110010000100110", 
	 "0110010000011110", 
	 "0110010000010110", 
	 "0110010000001111", 
	 "0110010000000111", 
	 "0110001111111111", 
	 "0110001111110111", 
	 "0110001111101111", 
	 "0110001111100111", 
	 "0110001111011111", 
	 "0110001111011000", 
	 "0110001111010000", 
	 "0110001111001000", 
	 "0110001111000000", 
	 "0110001110111000", 
	 "0110001110110000", 
	 "0110001110101000", 
	 "0110001110100000", 
	 "0110001110011001", 
	 "0110001110010001", 
	 "0110001110001001", 
	 "0110001110000001", 
	 "0110001101111001", 
	 "0110001101110001", 
	 "0110001101101001", 
	 "0110001101100001", 
	 "0110001101011001", 
	 "0110001101010001", 
	 "0110001101001001", 
	 "0110001101000010", 
	 "0110001100111010", 
	 "0110001100110010", 
	 "0110001100101010", 
	 "0110001100100010", 
	 "0110001100011010", 
	 "0110001100010010", 
	 "0110001100001010", 
	 "0110001100000010", 
	 "0110001011111010", 
	 "0110001011110010", 
	 "0110001011101010", 
	 "0110001011100010", 
	 "0110001011011010", 
	 "0110001011010010", 
	 "0110001011001010", 
	 "0110001011000010", 
	 "0110001010111010", 
	 "0110001010110010", 
	 "0110001010101010", 
	 "0110001010100010", 
	 "0110001010011010", 
	 "0110001010010010", 
	 "0110001010001010", 
	 "0110001010000010", 
	 "0110001001111010", 
	 "0110001001110010", 
	 "0110001001101010", 
	 "0110001001100010", 
	 "0110001001011010", 
	 "0110001001010010", 
	 "0110001001001010", 
	 "0110001001000010", 
	 "0110001000111010", 
	 "0110001000110010", 
	 "0110001000101010", 
	 "0110001000100001", 
	 "0110001000011001", 
	 "0110001000010001", 
	 "0110001000001001", 
	 "0110001000000001", 
	 "0110000111111001", 
	 "0110000111110001", 
	 "0110000111101001", 
	 "0110000111100001", 
	 "0110000111011001", 
	 "0110000111010001", 
	 "0110000111001001", 
	 "0110000111000000", 
	 "0110000110111000", 
	 "0110000110110000", 
	 "0110000110101000", 
	 "0110000110100000", 
	 "0110000110011000", 
	 "0110000110010000", 
	 "0110000110001000", 
	 "0110000101111111", 
	 "0110000101110111", 
	 "0110000101101111", 
	 "0110000101100111", 
	 "0110000101011111", 
	 "0110000101010111", 
	 "0110000101001110", 
	 "0110000101000110", 
	 "0110000100111110", 
	 "0110000100110110", 
	 "0110000100101110", 
	 "0110000100100110", 
	 "0110000100011101", 
	 "0110000100010101", 
	 "0110000100001101", 
	 "0110000100000101", 
	 "0110000011111101", 
	 "0110000011110100", 
	 "0110000011101100", 
	 "0110000011100100", 
	 "0110000011011100", 
	 "0110000011010100", 
	 "0110000011001011", 
	 "0110000011000011", 
	 "0110000010111011", 
	 "0110000010110011", 
	 "0110000010101010", 
	 "0110000010100010", 
	 "0110000010011010", 
	 "0110000010010010", 
	 "0110000010001001", 
	 "0110000010000001", 
	 "0110000001111001", 
	 "0110000001110001", 
	 "0110000001101000", 
	 "0110000001100000", 
	 "0110000001011000", 
	 "0110000001010000", 
	 "0110000001000111", 
	 "0110000000111111", 
	 "0110000000110111", 
	 "0110000000101110", 
	 "0110000000100110", 
	 "0110000000011110", 
	 "0110000000010110", 
	 "0110000000001101", 
	 "0110000000000101", 
	 "0101111111111101", 
	 "0101111111110100", 
	 "0101111111101100", 
	 "0101111111100100", 
	 "0101111111011011", 
	 "0101111111010011", 
	 "0101111111001011", 
	 "0101111111000010", 
	 "0101111110111010", 
	 "0101111110110010", 
	 "0101111110101001", 
	 "0101111110100001", 
	 "0101111110011001", 
	 "0101111110010000", 
	 "0101111110001000", 
	 "0101111110000000", 
	 "0101111101110111", 
	 "0101111101101111", 
	 "0101111101100110", 
	 "0101111101011110", 
	 "0101111101010110", 
	 "0101111101001101", 
	 "0101111101000101", 
	 "0101111100111100", 
	 "0101111100110100", 
	 "0101111100101100", 
	 "0101111100100011", 
	 "0101111100011011", 
	 "0101111100010010", 
	 "0101111100001010", 
	 "0101111100000010", 
	 "0101111011111001", 
	 "0101111011110001", 
	 "0101111011101000", 
	 "0101111011100000", 
	 "0101111011010111", 
	 "0101111011001111", 
	 "0101111011000111", 
	 "0101111010111110", 
	 "0101111010110110", 
	 "0101111010101101", 
	 "0101111010100101", 
	 "0101111010011100", 
	 "0101111010010100", 
	 "0101111010001011", 
	 "0101111010000011", 
	 "0101111001111010", 
	 "0101111001110010", 
	 "0101111001101001", 
	 "0101111001100001", 
	 "0101111001011000", 
	 "0101111001010000", 
	 "0101111001001000", 
	 "0101111000111111", 
	 "0101111000110111", 
	 "0101111000101110", 
	 "0101111000100101", 
	 "0101111000011101", 
	 "0101111000010100", 
	 "0101111000001100", 
	 "0101111000000011", 
	 "0101110111111011", 
	 "0101110111110010", 
	 "0101110111101010", 
	 "0101110111100001", 
	 "0101110111011001", 
	 "0101110111010000", 
	 "0101110111001000", 
	 "0101110110111111", 
	 "0101110110110111", 
	 "0101110110101110", 
	 "0101110110100101", 
	 "0101110110011101", 
	 "0101110110010100", 
	 "0101110110001100", 
	 "0101110110000011", 
	 "0101110101111010", 
	 "0101110101110010", 
	 "0101110101101001", 
	 "0101110101100001", 
	 "0101110101011000", 
	 "0101110101010000", 
	 "0101110101000111", 
	 "0101110100111110", 
	 "0101110100110110", 
	 "0101110100101101", 
	 "0101110100100100", 
	 "0101110100011100", 
	 "0101110100010011", 
	 "0101110100001011", 
	 "0101110100000010", 
	 "0101110011111001", 
	 "0101110011110001", 
	 "0101110011101000", 
	 "0101110011011111", 
	 "0101110011010111", 
	 "0101110011001110", 
	 "0101110011000101", 
	 "0101110010111101", 
	 "0101110010110100", 
	 "0101110010101011", 
	 "0101110010100011", 
	 "0101110010011010", 
	 "0101110010010001", 
	 "0101110010001001", 
	 "0101110010000000", 
	 "0101110001110111", 
	 "0101110001101111", 
	 "0101110001100110", 
	 "0101110001011101", 
	 "0101110001010101", 
	 "0101110001001100", 
	 "0101110001000011", 
	 "0101110000111010", 
	 "0101110000110010", 
	 "0101110000101001", 
	 "0101110000100000", 
	 "0101110000011000", 
	 "0101110000001111", 
	 "0101110000000110", 
	 "0101101111111101", 
	 "0101101111110101", 
	 "0101101111101100", 
	 "0101101111100011", 
	 "0101101111011010", 
	 "0101101111010010", 
	 "0101101111001001", 
	 "0101101111000000", 
	 "0101101110110111", 
	 "0101101110101111", 
	 "0101101110100110", 
	 "0101101110011101", 
	 "0101101110010100", 
	 "0101101110001100", 
	 "0101101110000011", 
	 "0101101101111010", 
	 "0101101101110001", 
	 "0101101101101000", 
	 "0101101101100000", 
	 "0101101101010111", 
	 "0101101101001110", 
	 "0101101101000101", 
	 "0101101100111100", 
	 "0101101100110100", 
	 "0101101100101011", 
	 "0101101100100010", 
	 "0101101100011001", 
	 "0101101100010000", 
	 "0101101100000111", 
	 "0101101011111111", 
	 "0101101011110110", 
	 "0101101011101101", 
	 "0101101011100100", 
	 "0101101011011011", 
	 "0101101011010010", 
	 "0101101011001001", 
	 "0101101011000001", 
	 "0101101010111000", 
	 "0101101010101111", 
	 "0101101010100110", 
	 "0101101010011101", 
	 "0101101010010100", 
	 "0101101010001011", 
	 "0101101010000010", 
	 "0101101001111010", 
	 "0101101001110001", 
	 "0101101001101000", 
	 "0101101001011111", 
	 "0101101001010110", 
	 "0101101001001101", 
	 "0101101001000100", 
	 "0101101000111011", 
	 "0101101000110010", 
	 "0101101000101001", 
	 "0101101000100001", 
	 "0101101000011000", 
	 "0101101000001111", 
	 "0101101000000110", 
	 "0101100111111101", 
	 "0101100111110100", 
	 "0101100111101011", 
	 "0101100111100010", 
	 "0101100111011001", 
	 "0101100111010000", 
	 "0101100111000111", 
	 "0101100110111110", 
	 "0101100110110101", 
	 "0101100110101100", 
	 "0101100110100011", 
	 "0101100110011010", 
	 "0101100110010001", 
	 "0101100110001000", 
	 "0101100101111111", 
	 "0101100101110110", 
	 "0101100101101101", 
	 "0101100101100100", 
	 "0101100101011011", 
	 "0101100101010010", 
	 "0101100101001001", 
	 "0101100101000000", 
	 "0101100100110111", 
	 "0101100100101110", 
	 "0101100100100101", 
	 "0101100100011100", 
	 "0101100100010011", 
	 "0101100100001010", 
	 "0101100100000001", 
	 "0101100011111000", 
	 "0101100011101111", 
	 "0101100011100110", 
	 "0101100011011101", 
	 "0101100011010100", 
	 "0101100011001011", 
	 "0101100011000010", 
	 "0101100010111001", 
	 "0101100010110000", 
	 "0101100010100111", 
	 "0101100010011110", 
	 "0101100010010101", 
	 "0101100010001100", 
	 "0101100010000010", 
	 "0101100001111001", 
	 "0101100001110000", 
	 "0101100001100111", 
	 "0101100001011110", 
	 "0101100001010101", 
	 "0101100001001100", 
	 "0101100001000011", 
	 "0101100000111010", 
	 "0101100000110001", 
	 "0101100000101000", 
	 "0101100000011110", 
	 "0101100000010101", 
	 "0101100000001100", 
	 "0101100000000011", 
	 "0101011111111010", 
	 "0101011111110001", 
	 "0101011111101000", 
	 "0101011111011111", 
	 "0101011111010101", 
	 "0101011111001100", 
	 "0101011111000011", 
	 "0101011110111010", 
	 "0101011110110001", 
	 "0101011110101000", 
	 "0101011110011111", 
	 "0101011110010101", 
	 "0101011110001100", 
	 "0101011110000011", 
	 "0101011101111010", 
	 "0101011101110001", 
	 "0101011101100111", 
	 "0101011101011110", 
	 "0101011101010101", 
	 "0101011101001100", 
	 "0101011101000011", 
	 "0101011100111010", 
	 "0101011100110000", 
	 "0101011100100111", 
	 "0101011100011110", 
	 "0101011100010101", 
	 "0101011100001100", 
	 "0101011100000010", 
	 "0101011011111001", 
	 "0101011011110000", 
	 "0101011011100111", 
	 "0101011011011101", 
	 "0101011011010100", 
	 "0101011011001011", 
	 "0101011011000010", 
	 "0101011010111000", 
	 "0101011010101111", 
	 "0101011010100110", 
	 "0101011010011101", 
	 "0101011010010011", 
	 "0101011010001010", 
	 "0101011010000001", 
	 "0101011001111000", 
	 "0101011001101110", 
	 "0101011001100101", 
	 "0101011001011100", 
	 "0101011001010011", 
	 "0101011001001001", 
	 "0101011001000000", 
	 "0101011000110111", 
	 "0101011000101101", 
	 "0101011000100100", 
	 "0101011000011011", 
	 "0101011000010010", 
	 "0101011000001000", 
	 "0101010111111111", 
	 "0101010111110110", 
	 "0101010111101100", 
	 "0101010111100011", 
	 "0101010111011010", 
	 "0101010111010000", 
	 "0101010111000111", 
	 "0101010110111110", 
	 "0101010110110100", 
	 "0101010110101011", 
	 "0101010110100010", 
	 "0101010110011000", 
	 "0101010110001111", 
	 "0101010110000110", 
	 "0101010101111100", 
	 "0101010101110011", 
	 "0101010101101010", 
	 "0101010101100000", 
	 "0101010101010111", 
	 "0101010101001110", 
	 "0101010101000100", 
	 "0101010100111011", 
	 "0101010100110001", 
	 "0101010100101000", 
	 "0101010100011111", 
	 "0101010100010101", 
	 "0101010100001100", 
	 "0101010100000010", 
	 "0101010011111001", 
	 "0101010011110000", 
	 "0101010011100110", 
	 "0101010011011101", 
	 "0101010011010011", 
	 "0101010011001010", 
	 "0101010011000001", 
	 "0101010010110111", 
	 "0101010010101110", 
	 "0101010010100100", 
	 "0101010010011011", 
	 "0101010010010001", 
	 "0101010010001000", 
	 "0101010001111111", 
	 "0101010001110101", 
	 "0101010001101100", 
	 "0101010001100010", 
	 "0101010001011001", 
	 "0101010001001111", 
	 "0101010001000110", 
	 "0101010000111100", 
	 "0101010000110011", 
	 "0101010000101010", 
	 "0101010000100000", 
	 "0101010000010111", 
	 "0101010000001101", 
	 "0101010000000100", 
	 "0101001111111010", 
	 "0101001111110001", 
	 "0101001111100111", 
	 "0101001111011110", 
	 "0101001111010100", 
	 "0101001111001011", 
	 "0101001111000001", 
	 "0101001110111000", 
	 "0101001110101110", 
	 "0101001110100101", 
	 "0101001110011011", 
	 "0101001110010010", 
	 "0101001110001000", 
	 "0101001101111111", 
	 "0101001101110101", 
	 "0101001101101100", 
	 "0101001101100010", 
	 "0101001101011000", 
	 "0101001101001111", 
	 "0101001101000101", 
	 "0101001100111100", 
	 "0101001100110010", 
	 "0101001100101001", 
	 "0101001100011111", 
	 "0101001100010110", 
	 "0101001100001100", 
	 "0101001100000011", 
	 "0101001011111001", 
	 "0101001011101111", 
	 "0101001011100110", 
	 "0101001011011100", 
	 "0101001011010011", 
	 "0101001011001001", 
	 "0101001010111111", 
	 "0101001010110110", 
	 "0101001010101100", 
	 "0101001010100011", 
	 "0101001010011001", 
	 "0101001010010000", 
	 "0101001010000110", 
	 "0101001001111100", 
	 "0101001001110011", 
	 "0101001001101001", 
	 "0101001001011111", 
	 "0101001001010110", 
	 "0101001001001100", 
	 "0101001001000011", 
	 "0101001000111001", 
	 "0101001000101111", 
	 "0101001000100110", 
	 "0101001000011100", 
	 "0101001000010010", 
	 "0101001000001001", 
	 "0101000111111111", 
	 "0101000111110101", 
	 "0101000111101100", 
	 "0101000111100010", 
	 "0101000111011000", 
	 "0101000111001111", 
	 "0101000111000101", 
	 "0101000110111011", 
	 "0101000110110010", 
	 "0101000110101000", 
	 "0101000110011110", 
	 "0101000110010101", 
	 "0101000110001011", 
	 "0101000110000001", 
	 "0101000101111000", 
	 "0101000101101110", 
	 "0101000101100100", 
	 "0101000101011011", 
	 "0101000101010001", 
	 "0101000101000111", 
	 "0101000100111110", 
	 "0101000100110100", 
	 "0101000100101010", 
	 "0101000100100000", 
	 "0101000100010111", 
	 "0101000100001101", 
	 "0101000100000011", 
	 "0101000011111001", 
	 "0101000011110000", 
	 "0101000011100110", 
	 "0101000011011100", 
	 "0101000011010011", 
	 "0101000011001001", 
	 "0101000010111111", 
	 "0101000010110101", 
	 "0101000010101100", 
	 "0101000010100010", 
	 "0101000010011000", 
	 "0101000010001110", 
	 "0101000010000100", 
	 "0101000001111011", 
	 "0101000001110001", 
	 "0101000001100111", 
	 "0101000001011101", 
	 "0101000001010100", 
	 "0101000001001010", 
	 "0101000001000000", 
	 "0101000000110110", 
	 "0101000000101100", 
	 "0101000000100011", 
	 "0101000000011001", 
	 "0101000000001111", 
	 "0101000000000101", 
	 "0100111111111011", 
	 "0100111111110010", 
	 "0100111111101000", 
	 "0100111111011110", 
	 "0100111111010100", 
	 "0100111111001010", 
	 "0100111111000000", 
	 "0100111110110111", 
	 "0100111110101101", 
	 "0100111110100011", 
	 "0100111110011001", 
	 "0100111110001111", 
	 "0100111110000101", 
	 "0100111101111100", 
	 "0100111101110010", 
	 "0100111101101000", 
	 "0100111101011110", 
	 "0100111101010100", 
	 "0100111101001010", 
	 "0100111101000000", 
	 "0100111100110111", 
	 "0100111100101101", 
	 "0100111100100011", 
	 "0100111100011001", 
	 "0100111100001111", 
	 "0100111100000101", 
	 "0100111011111011", 
	 "0100111011110001", 
	 "0100111011101000", 
	 "0100111011011110", 
	 "0100111011010100", 
	 "0100111011001010", 
	 "0100111011000000", 
	 "0100111010110110", 
	 "0100111010101100", 
	 "0100111010100010", 
	 "0100111010011000", 
	 "0100111010001110", 
	 "0100111010000100", 
	 "0100111001111010", 
	 "0100111001110001", 
	 "0100111001100111", 
	 "0100111001011101", 
	 "0100111001010011", 
	 "0100111001001001", 
	 "0100111000111111", 
	 "0100111000110101", 
	 "0100111000101011", 
	 "0100111000100001", 
	 "0100111000010111", 
	 "0100111000001101", 
	 "0100111000000011", 
	 "0100110111111001", 
	 "0100110111101111", 
	 "0100110111100101", 
	 "0100110111011011", 
	 "0100110111010001", 
	 "0100110111000111", 
	 "0100110110111101", 
	 "0100110110110011", 
	 "0100110110101001", 
	 "0100110110011111", 
	 "0100110110010101", 
	 "0100110110001011", 
	 "0100110110000001", 
	 "0100110101110111", 
	 "0100110101101101", 
	 "0100110101100011", 
	 "0100110101011001", 
	 "0100110101001111", 
	 "0100110101000101", 
	 "0100110100111011", 
	 "0100110100110001", 
	 "0100110100100111", 
	 "0100110100011101", 
	 "0100110100010011", 
	 "0100110100001001", 
	 "0100110011111111", 
	 "0100110011110101", 
	 "0100110011101011", 
	 "0100110011100001", 
	 "0100110011010111", 
	 "0100110011001101", 
	 "0100110011000011", 
	 "0100110010111001", 
	 "0100110010101111", 
	 "0100110010100101", 
	 "0100110010011011", 
	 "0100110010010001", 
	 "0100110010000110", 
	 "0100110001111100", 
	 "0100110001110010", 
	 "0100110001101000", 
	 "0100110001011110", 
	 "0100110001010100", 
	 "0100110001001010", 
	 "0100110001000000", 
	 "0100110000110110", 
	 "0100110000101100", 
	 "0100110000100010", 
	 "0100110000010111", 
	 "0100110000001101", 
	 "0100110000000011", 
	 "0100101111111001", 
	 "0100101111101111", 
	 "0100101111100101", 
	 "0100101111011011", 
	 "0100101111010001", 
	 "0100101111000111", 
	 "0100101110111100", 
	 "0100101110110010", 
	 "0100101110101000", 
	 "0100101110011110", 
	 "0100101110010100", 
	 "0100101110001010", 
	 "0100101110000000", 
	 "0100101101110101", 
	 "0100101101101011", 
	 "0100101101100001", 
	 "0100101101010111", 
	 "0100101101001101", 
	 "0100101101000011", 
	 "0100101100111000", 
	 "0100101100101110", 
	 "0100101100100100", 
	 "0100101100011010", 
	 "0100101100010000", 
	 "0100101100000110", 
	 "0100101011111011", 
	 "0100101011110001", 
	 "0100101011100111", 
	 "0100101011011101", 
	 "0100101011010011", 
	 "0100101011001000", 
	 "0100101010111110", 
	 "0100101010110100", 
	 "0100101010101010", 
	 "0100101010100000", 
	 "0100101010010101", 
	 "0100101010001011", 
	 "0100101010000001", 
	 "0100101001110111", 
	 "0100101001101101", 
	 "0100101001100010", 
	 "0100101001011000", 
	 "0100101001001110", 
	 "0100101001000100", 
	 "0100101000111001", 
	 "0100101000101111", 
	 "0100101000100101", 
	 "0100101000011011", 
	 "0100101000010000", 
	 "0100101000000110", 
	 "0100100111111100", 
	 "0100100111110010", 
	 "0100100111100111", 
	 "0100100111011101", 
	 "0100100111010011", 
	 "0100100111001001", 
	 "0100100110111110", 
	 "0100100110110100", 
	 "0100100110101010", 
	 "0100100110100000", 
	 "0100100110010101", 
	 "0100100110001011", 
	 "0100100110000001", 
	 "0100100101110110", 
	 "0100100101101100", 
	 "0100100101100010", 
	 "0100100101011000", 
	 "0100100101001101", 
	 "0100100101000011", 
	 "0100100100111001", 
	 "0100100100101110", 
	 "0100100100100100", 
	 "0100100100011010", 
	 "0100100100001111", 
	 "0100100100000101", 
	 "0100100011111011", 
	 "0100100011110000", 
	 "0100100011100110", 
	 "0100100011011100", 
	 "0100100011010001", 
	 "0100100011000111", 
	 "0100100010111101", 
	 "0100100010110010", 
	 "0100100010101000", 
	 "0100100010011110", 
	 "0100100010010011", 
	 "0100100010001001", 
	 "0100100001111111", 
	 "0100100001110100", 
	 "0100100001101010", 
	 "0100100001100000", 
	 "0100100001010101", 
	 "0100100001001011", 
	 "0100100001000000", 
	 "0100100000110110", 
	 "0100100000101100", 
	 "0100100000100001", 
	 "0100100000010111", 
	 "0100100000001101", 
	 "0100100000000010", 
	 "0100011111111000", 
	 "0100011111101101", 
	 "0100011111100011", 
	 "0100011111011001", 
	 "0100011111001110", 
	 "0100011111000100", 
	 "0100011110111001", 
	 "0100011110101111", 
	 "0100011110100101", 
	 "0100011110011010", 
	 "0100011110010000", 
	 "0100011110000101", 
	 "0100011101111011", 
	 "0100011101110000", 
	 "0100011101100110", 
	 "0100011101011100", 
	 "0100011101010001", 
	 "0100011101000111", 
	 "0100011100111100", 
	 "0100011100110010", 
	 "0100011100100111", 
	 "0100011100011101", 
	 "0100011100010010", 
	 "0100011100001000", 
	 "0100011011111110", 
	 "0100011011110011", 
	 "0100011011101001", 
	 "0100011011011110", 
	 "0100011011010100", 
	 "0100011011001001", 
	 "0100011010111111", 
	 "0100011010110100", 
	 "0100011010101010", 
	 "0100011010011111", 
	 "0100011010010101", 
	 "0100011010001010", 
	 "0100011010000000", 
	 "0100011001110101", 
	 "0100011001101011", 
	 "0100011001100000", 
	 "0100011001010110", 
	 "0100011001001011", 
	 "0100011001000001", 
	 "0100011000110110", 
	 "0100011000101100", 
	 "0100011000100001", 
	 "0100011000010111", 
	 "0100011000001100", 
	 "0100011000000010", 
	 "0100010111110111", 
	 "0100010111101101", 
	 "0100010111100010", 
	 "0100010111011000", 
	 "0100010111001101", 
	 "0100010111000011", 
	 "0100010110111000", 
	 "0100010110101110", 
	 "0100010110100011", 
	 "0100010110011001", 
	 "0100010110001110", 
	 "0100010110000011", 
	 "0100010101111001", 
	 "0100010101101110", 
	 "0100010101100100", 
	 "0100010101011001", 
	 "0100010101001111", 
	 "0100010101000100", 
	 "0100010100111001", 
	 "0100010100101111", 
	 "0100010100100100", 
	 "0100010100011010", 
	 "0100010100001111", 
	 "0100010100000101", 
	 "0100010011111010", 
	 "0100010011101111", 
	 "0100010011100101", 
	 "0100010011011010", 
	 "0100010011010000", 
	 "0100010011000101", 
	 "0100010010111010", 
	 "0100010010110000", 
	 "0100010010100101", 
	 "0100010010011011", 
	 "0100010010010000", 
	 "0100010010000101", 
	 "0100010001111011", 
	 "0100010001110000", 
	 "0100010001100110", 
	 "0100010001011011", 
	 "0100010001010000", 
	 "0100010001000110", 
	 "0100010000111011", 
	 "0100010000110000", 
	 "0100010000100110", 
	 "0100010000011011", 
	 "0100010000010001", 
	 "0100010000000110", 
	 "0100001111111011", 
	 "0100001111110001", 
	 "0100001111100110", 
	 "0100001111011011", 
	 "0100001111010001", 
	 "0100001111000110", 
	 "0100001110111011", 
	 "0100001110110001", 
	 "0100001110100110", 
	 "0100001110011011", 
	 "0100001110010001", 
	 "0100001110000110", 
	 "0100001101111011", 
	 "0100001101110001", 
	 "0100001101100110", 
	 "0100001101011011", 
	 "0100001101010001", 
	 "0100001101000110", 
	 "0100001100111011", 
	 "0100001100110000", 
	 "0100001100100110", 
	 "0100001100011011", 
	 "0100001100010000", 
	 "0100001100000110", 
	 "0100001011111011", 
	 "0100001011110000", 
	 "0100001011100110", 
	 "0100001011011011", 
	 "0100001011010000", 
	 "0100001011000101", 
	 "0100001010111011", 
	 "0100001010110000", 
	 "0100001010100101", 
	 "0100001010011010", 
	 "0100001010010000", 
	 "0100001010000101", 
	 "0100001001111010", 
	 "0100001001110000", 
	 "0100001001100101", 
	 "0100001001011010", 
	 "0100001001001111", 
	 "0100001001000101", 
	 "0100001000111010", 
	 "0100001000101111", 
	 "0100001000100100", 
	 "0100001000011010", 
	 "0100001000001111", 
	 "0100001000000100", 
	 "0100000111111001", 
	 "0100000111101110", 
	 "0100000111100100", 
	 "0100000111011001", 
	 "0100000111001110", 
	 "0100000111000011", 
	 "0100000110111001", 
	 "0100000110101110", 
	 "0100000110100011", 
	 "0100000110011000", 
	 "0100000110001101", 
	 "0100000110000011", 
	 "0100000101111000", 
	 "0100000101101101", 
	 "0100000101100010", 
	 "0100000101010111", 
	 "0100000101001101", 
	 "0100000101000010", 
	 "0100000100110111", 
	 "0100000100101100", 
	 "0100000100100001", 
	 "0100000100010111", 
	 "0100000100001100", 
	 "0100000100000001", 
	 "0100000011110110", 
	 "0100000011101011", 
	 "0100000011100000", 
	 "0100000011010110", 
	 "0100000011001011", 
	 "0100000011000000", 
	 "0100000010110101", 
	 "0100000010101010", 
	 "0100000010011111", 
	 "0100000010010101", 
	 "0100000010001010", 
	 "0100000001111111", 
	 "0100000001110100", 
	 "0100000001101001", 
	 "0100000001011110", 
	 "0100000001010011", 
	 "0100000001001000", 
	 "0100000000111110", 
	 "0100000000110011", 
	 "0100000000101000", 
	 "0100000000011101", 
	 "0100000000010010", 
	 "0100000000000111", 
	 "0011111111111100", 
	 "0011111111110001", 
	 "0011111111100111", 
	 "0011111111011100", 
	 "0011111111010001", 
	 "0011111111000110", 
	 "0011111110111011", 
	 "0011111110110000", 
	 "0011111110100101", 
	 "0011111110011010", 
	 "0011111110001111", 
	 "0011111110000101", 
	 "0011111101111010", 
	 "0011111101101111", 
	 "0011111101100100", 
	 "0011111101011001", 
	 "0011111101001110", 
	 "0011111101000011", 
	 "0011111100111000", 
	 "0011111100101101", 
	 "0011111100100010", 
	 "0011111100010111", 
	 "0011111100001100", 
	 "0011111100000001", 
	 "0011111011110110", 
	 "0011111011101100", 
	 "0011111011100001", 
	 "0011111011010110", 
	 "0011111011001011", 
	 "0011111011000000", 
	 "0011111010110101", 
	 "0011111010101010", 
	 "0011111010011111", 
	 "0011111010010100", 
	 "0011111010001001", 
	 "0011111001111110", 
	 "0011111001110011", 
	 "0011111001101000", 
	 "0011111001011101", 
	 "0011111001010010", 
	 "0011111001000111", 
	 "0011111000111100", 
	 "0011111000110001", 
	 "0011111000100110", 
	 "0011111000011011", 
	 "0011111000010000", 
	 "0011111000000101", 
	 "0011110111111010", 
	 "0011110111101111", 
	 "0011110111100100", 
	 "0011110111011001", 
	 "0011110111001110", 
	 "0011110111000011", 
	 "0011110110111000", 
	 "0011110110101101", 
	 "0011110110100010", 
	 "0011110110010111", 
	 "0011110110001100", 
	 "0011110110000001", 
	 "0011110101110110", 
	 "0011110101101011", 
	 "0011110101100000", 
	 "0011110101010101", 
	 "0011110101001010", 
	 "0011110100111111", 
	 "0011110100110100", 
	 "0011110100101001", 
	 "0011110100011110", 
	 "0011110100010011", 
	 "0011110100001000", 
	 "0011110011111101", 
	 "0011110011110010", 
	 "0011110011100111", 
	 "0011110011011100", 
	 "0011110011010000", 
	 "0011110011000101", 
	 "0011110010111010", 
	 "0011110010101111", 
	 "0011110010100100", 
	 "0011110010011001", 
	 "0011110010001110", 
	 "0011110010000011", 
	 "0011110001111000", 
	 "0011110001101101", 
	 "0011110001100010", 
	 "0011110001010111", 
	 "0011110001001100", 
	 "0011110001000001", 
	 "0011110000110101", 
	 "0011110000101010", 
	 "0011110000011111", 
	 "0011110000010100", 
	 "0011110000001001", 
	 "0011101111111110", 
	 "0011101111110011", 
	 "0011101111101000", 
	 "0011101111011101", 
	 "0011101111010010", 
	 "0011101111000110", 
	 "0011101110111011", 
	 "0011101110110000", 
	 "0011101110100101", 
	 "0011101110011010", 
	 "0011101110001111", 
	 "0011101110000100", 
	 "0011101101111001", 
	 "0011101101101101", 
	 "0011101101100010", 
	 "0011101101010111", 
	 "0011101101001100", 
	 "0011101101000001", 
	 "0011101100110110", 
	 "0011101100101011", 
	 "0011101100100000", 
	 "0011101100010100", 
	 "0011101100001001", 
	 "0011101011111110", 
	 "0011101011110011", 
	 "0011101011101000", 
	 "0011101011011101", 
	 "0011101011010001", 
	 "0011101011000110", 
	 "0011101010111011", 
	 "0011101010110000", 
	 "0011101010100101", 
	 "0011101010011010", 
	 "0011101010001110", 
	 "0011101010000011", 
	 "0011101001111000", 
	 "0011101001101101", 
	 "0011101001100010", 
	 "0011101001010111", 
	 "0011101001001011", 
	 "0011101001000000", 
	 "0011101000110101", 
	 "0011101000101010", 
	 "0011101000011111", 
	 "0011101000010011", 
	 "0011101000001000", 
	 "0011100111111101", 
	 "0011100111110010", 
	 "0011100111100111", 
	 "0011100111011011", 
	 "0011100111010000", 
	 "0011100111000101", 
	 "0011100110111010", 
	 "0011100110101111", 
	 "0011100110100011", 
	 "0011100110011000", 
	 "0011100110001101", 
	 "0011100110000010", 
	 "0011100101110110", 
	 "0011100101101011", 
	 "0011100101100000", 
	 "0011100101010101", 
	 "0011100101001001", 
	 "0011100100111110", 
	 "0011100100110011", 
	 "0011100100101000", 
	 "0011100100011101", 
	 "0011100100010001", 
	 "0011100100000110", 
	 "0011100011111011", 
	 "0011100011110000", 
	 "0011100011100100", 
	 "0011100011011001", 
	 "0011100011001110", 
	 "0011100011000010", 
	 "0011100010110111", 
	 "0011100010101100", 
	 "0011100010100001", 
	 "0011100010010101", 
	 "0011100010001010", 
	 "0011100001111111", 
	 "0011100001110100", 
	 "0011100001101000", 
	 "0011100001011101", 
	 "0011100001010010", 
	 "0011100001000110", 
	 "0011100000111011", 
	 "0011100000110000", 
	 "0011100000100101", 
	 "0011100000011001", 
	 "0011100000001110", 
	 "0011100000000011", 
	 "0011011111110111", 
	 "0011011111101100", 
	 "0011011111100001", 
	 "0011011111010101", 
	 "0011011111001010", 
	 "0011011110111111", 
	 "0011011110110100", 
	 "0011011110101000", 
	 "0011011110011101", 
	 "0011011110010010", 
	 "0011011110000110", 
	 "0011011101111011", 
	 "0011011101110000", 
	 "0011011101100100", 
	 "0011011101011001", 
	 "0011011101001110", 
	 "0011011101000010", 
	 "0011011100110111", 
	 "0011011100101100", 
	 "0011011100100000", 
	 "0011011100010101", 
	 "0011011100001010", 
	 "0011011011111110", 
	 "0011011011110011", 
	 "0011011011101000", 
	 "0011011011011100", 
	 "0011011011010001", 
	 "0011011011000101", 
	 "0011011010111010", 
	 "0011011010101111", 
	 "0011011010100011", 
	 "0011011010011000", 
	 "0011011010001101", 
	 "0011011010000001", 
	 "0011011001110110", 
	 "0011011001101011", 
	 "0011011001011111", 
	 "0011011001010100", 
	 "0011011001001000", 
	 "0011011000111101", 
	 "0011011000110010", 
	 "0011011000100110", 
	 "0011011000011011", 
	 "0011011000001111", 
	 "0011011000000100", 
	 "0011010111111001", 
	 "0011010111101101", 
	 "0011010111100010", 
	 "0011010111010111", 
	 "0011010111001011", 
	 "0011010111000000", 
	 "0011010110110100", 
	 "0011010110101001", 
	 "0011010110011101", 
	 "0011010110010010", 
	 "0011010110000111", 
	 "0011010101111011", 
	 "0011010101110000", 
	 "0011010101100100", 
	 "0011010101011001", 
	 "0011010101001110", 
	 "0011010101000010", 
	 "0011010100110111", 
	 "0011010100101011", 
	 "0011010100100000", 
	 "0011010100010100", 
	 "0011010100001001", 
	 "0011010011111110", 
	 "0011010011110010", 
	 "0011010011100111", 
	 "0011010011011011", 
	 "0011010011010000", 
	 "0011010011000100", 
	 "0011010010111001", 
	 "0011010010101101", 
	 "0011010010100010", 
	 "0011010010010111", 
	 "0011010010001011", 
	 "0011010010000000", 
	 "0011010001110100", 
	 "0011010001101001", 
	 "0011010001011101", 
	 "0011010001010010", 
	 "0011010001000110", 
	 "0011010000111011", 
	 "0011010000101111", 
	 "0011010000100100", 
	 "0011010000011000", 
	 "0011010000001101", 
	 "0011010000000001", 
	 "0011001111110110", 
	 "0011001111101010", 
	 "0011001111011111", 
	 "0011001111010011", 
	 "0011001111001000", 
	 "0011001110111100", 
	 "0011001110110001", 
	 "0011001110100101", 
	 "0011001110011010", 
	 "0011001110001110", 
	 "0011001110000011", 
	 "0011001101110111", 
	 "0011001101101100", 
	 "0011001101100000", 
	 "0011001101010101", 
	 "0011001101001001", 
	 "0011001100111110", 
	 "0011001100110010", 
	 "0011001100100111", 
	 "0011001100011011", 
	 "0011001100010000", 
	 "0011001100000100", 
	 "0011001011111001", 
	 "0011001011101101", 
	 "0011001011100010", 
	 "0011001011010110", 
	 "0011001011001011", 
	 "0011001010111111", 
	 "0011001010110100", 
	 "0011001010101000", 
	 "0011001010011101", 
	 "0011001010010001", 
	 "0011001010000101", 
	 "0011001001111010", 
	 "0011001001101110", 
	 "0011001001100011", 
	 "0011001001010111", 
	 "0011001001001100", 
	 "0011001001000000", 
	 "0011001000110101", 
	 "0011001000101001", 
	 "0011001000011101", 
	 "0011001000010010", 
	 "0011001000000110", 
	 "0011000111111011", 
	 "0011000111101111", 
	 "0011000111100100", 
	 "0011000111011000", 
	 "0011000111001100", 
	 "0011000111000001", 
	 "0011000110110101", 
	 "0011000110101010", 
	 "0011000110011110", 
	 "0011000110010011", 
	 "0011000110000111", 
	 "0011000101111011", 
	 "0011000101110000", 
	 "0011000101100100", 
	 "0011000101011001", 
	 "0011000101001101", 
	 "0011000101000001", 
	 "0011000100110110", 
	 "0011000100101010", 
	 "0011000100011111", 
	 "0011000100010011", 
	 "0011000100000111", 
	 "0011000011111100", 
	 "0011000011110000", 
	 "0011000011100101", 
	 "0011000011011001", 
	 "0011000011001101", 
	 "0011000011000010", 
	 "0011000010110110", 
	 "0011000010101010", 
	 "0011000010011111", 
	 "0011000010010011", 
	 "0011000010001000", 
	 "0011000001111100", 
	 "0011000001110000", 
	 "0011000001100101", 
	 "0011000001011001", 
	 "0011000001001101", 
	 "0011000001000010", 
	 "0011000000110110", 
	 "0011000000101010", 
	 "0011000000011111", 
	 "0011000000010011", 
	 "0011000000001000", 
	 "0010111111111100", 
	 "0010111111110000", 
	 "0010111111100101", 
	 "0010111111011001", 
	 "0010111111001101", 
	 "0010111111000010", 
	 "0010111110110110", 
	 "0010111110101010", 
	 "0010111110011111", 
	 "0010111110010011", 
	 "0010111110000111", 
	 "0010111101111100", 
	 "0010111101110000", 
	 "0010111101100100", 
	 "0010111101011001", 
	 "0010111101001101", 
	 "0010111101000001", 
	 "0010111100110110", 
	 "0010111100101010", 
	 "0010111100011110", 
	 "0010111100010011", 
	 "0010111100000111", 
	 "0010111011111011", 
	 "0010111011101111", 
	 "0010111011100100", 
	 "0010111011011000", 
	 "0010111011001100", 
	 "0010111011000001", 
	 "0010111010110101", 
	 "0010111010101001", 
	 "0010111010011110", 
	 "0010111010010010", 
	 "0010111010000110", 
	 "0010111001111010", 
	 "0010111001101111", 
	 "0010111001100011", 
	 "0010111001010111", 
	 "0010111001001100", 
	 "0010111001000000", 
	 "0010111000110100", 
	 "0010111000101000", 
	 "0010111000011101", 
	 "0010111000010001", 
	 "0010111000000101", 
	 "0010110111111010", 
	 "0010110111101110", 
	 "0010110111100010", 
	 "0010110111010110", 
	 "0010110111001011", 
	 "0010110110111111", 
	 "0010110110110011", 
	 "0010110110100111", 
	 "0010110110011100", 
	 "0010110110010000", 
	 "0010110110000100", 
	 "0010110101111000", 
	 "0010110101101101", 
	 "0010110101100001", 
	 "0010110101010101", 
	 "0010110101001001", 
	 "0010110100111110", 
	 "0010110100110010", 
	 "0010110100100110", 
	 "0010110100011010", 
	 "0010110100001111", 
	 "0010110100000011", 
	 "0010110011110111", 
	 "0010110011101011", 
	 "0010110011100000", 
	 "0010110011010100", 
	 "0010110011001000", 
	 "0010110010111100", 
	 "0010110010110001", 
	 "0010110010100101", 
	 "0010110010011001", 
	 "0010110010001101", 
	 "0010110010000001", 
	 "0010110001110110", 
	 "0010110001101010", 
	 "0010110001011110", 
	 "0010110001010010", 
	 "0010110001000110", 
	 "0010110000111011", 
	 "0010110000101111", 
	 "0010110000100011", 
	 "0010110000010111", 
	 "0010110000001100", 
	 "0010110000000000", 
	 "0010101111110100", 
	 "0010101111101000", 
	 "0010101111011100", 
	 "0010101111010000", 
	 "0010101111000101", 
	 "0010101110111001", 
	 "0010101110101101", 
	 "0010101110100001", 
	 "0010101110010101", 
	 "0010101110001010", 
	 "0010101101111110", 
	 "0010101101110010", 
	 "0010101101100110", 
	 "0010101101011010", 
	 "0010101101001111", 
	 "0010101101000011", 
	 "0010101100110111", 
	 "0010101100101011", 
	 "0010101100011111", 
	 "0010101100010011", 
	 "0010101100001000", 
	 "0010101011111100", 
	 "0010101011110000", 
	 "0010101011100100", 
	 "0010101011011000", 
	 "0010101011001100", 
	 "0010101011000001", 
	 "0010101010110101", 
	 "0010101010101001", 
	 "0010101010011101", 
	 "0010101010010001", 
	 "0010101010000101", 
	 "0010101001111001", 
	 "0010101001101110", 
	 "0010101001100010", 
	 "0010101001010110", 
	 "0010101001001010", 
	 "0010101000111110", 
	 "0010101000110010", 
	 "0010101000100110", 
	 "0010101000011011", 
	 "0010101000001111", 
	 "0010101000000011", 
	 "0010100111110111", 
	 "0010100111101011", 
	 "0010100111011111", 
	 "0010100111010011", 
	 "0010100111000111", 
	 "0010100110111100", 
	 "0010100110110000", 
	 "0010100110100100", 
	 "0010100110011000", 
	 "0010100110001100", 
	 "0010100110000000", 
	 "0010100101110100", 
	 "0010100101101000", 
	 "0010100101011100", 
	 "0010100101010001", 
	 "0010100101000101", 
	 "0010100100111001", 
	 "0010100100101101", 
	 "0010100100100001", 
	 "0010100100010101", 
	 "0010100100001001", 
	 "0010100011111101", 
	 "0010100011110001", 
	 "0010100011100101", 
	 "0010100011011010", 
	 "0010100011001110", 
	 "0010100011000010", 
	 "0010100010110110", 
	 "0010100010101010", 
	 "0010100010011110", 
	 "0010100010010010", 
	 "0010100010000110", 
	 "0010100001111010", 
	 "0010100001101110", 
	 "0010100001100010", 
	 "0010100001010110", 
	 "0010100001001011", 
	 "0010100000111111", 
	 "0010100000110011", 
	 "0010100000100111", 
	 "0010100000011011", 
	 "0010100000001111", 
	 "0010100000000011", 
	 "0010011111110111", 
	 "0010011111101011", 
	 "0010011111011111", 
	 "0010011111010011", 
	 "0010011111000111", 
	 "0010011110111011", 
	 "0010011110101111", 
	 "0010011110100011", 
	 "0010011110010111", 
	 "0010011110001011", 
	 "0010011110000000", 
	 "0010011101110100", 
	 "0010011101101000", 
	 "0010011101011100", 
	 "0010011101010000", 
	 "0010011101000100", 
	 "0010011100111000", 
	 "0010011100101100", 
	 "0010011100100000", 
	 "0010011100010100", 
	 "0010011100001000", 
	 "0010011011111100", 
	 "0010011011110000", 
	 "0010011011100100", 
	 "0010011011011000", 
	 "0010011011001100", 
	 "0010011011000000", 
	 "0010011010110100", 
	 "0010011010101000", 
	 "0010011010011100", 
	 "0010011010010000", 
	 "0010011010000100", 
	 "0010011001111000", 
	 "0010011001101100", 
	 "0010011001100000", 
	 "0010011001010100", 
	 "0010011001001000", 
	 "0010011000111100", 
	 "0010011000110000", 
	 "0010011000100100", 
	 "0010011000011000", 
	 "0010011000001100", 
	 "0010011000000000", 
	 "0010010111110100", 
	 "0010010111101000", 
	 "0010010111011100", 
	 "0010010111010000", 
	 "0010010111000100", 
	 "0010010110111000", 
	 "0010010110101100", 
	 "0010010110100000", 
	 "0010010110010100", 
	 "0010010110001000", 
	 "0010010101111100", 
	 "0010010101110000", 
	 "0010010101100100", 
	 "0010010101011000", 
	 "0010010101001100", 
	 "0010010101000000", 
	 "0010010100110100", 
	 "0010010100101000", 
	 "0010010100011100", 
	 "0010010100010000", 
	 "0010010100000100", 
	 "0010010011111000", 
	 "0010010011101100", 
	 "0010010011100000", 
	 "0010010011010100", 
	 "0010010011001000", 
	 "0010010010111100", 
	 "0010010010110000", 
	 "0010010010100100", 
	 "0010010010011000", 
	 "0010010010001100", 
	 "0010010010000000", 
	 "0010010001110100", 
	 "0010010001100111", 
	 "0010010001011011", 
	 "0010010001001111", 
	 "0010010001000011", 
	 "0010010000110111", 
	 "0010010000101011", 
	 "0010010000011111", 
	 "0010010000010011", 
	 "0010010000000111", 
	 "0010001111111011", 
	 "0010001111101111", 
	 "0010001111100011", 
	 "0010001111010111", 
	 "0010001111001011", 
	 "0010001110111111", 
	 "0010001110110011", 
	 "0010001110100111", 
	 "0010001110011010", 
	 "0010001110001110", 
	 "0010001110000010", 
	 "0010001101110110", 
	 "0010001101101010", 
	 "0010001101011110", 
	 "0010001101010010", 
	 "0010001101000110", 
	 "0010001100111010", 
	 "0010001100101110", 
	 "0010001100100010", 
	 "0010001100010110", 
	 "0010001100001010", 
	 "0010001011111101", 
	 "0010001011110001", 
	 "0010001011100101", 
	 "0010001011011001", 
	 "0010001011001101", 
	 "0010001011000001", 
	 "0010001010110101", 
	 "0010001010101001", 
	 "0010001010011101", 
	 "0010001010010001", 
	 "0010001010000100", 
	 "0010001001111000", 
	 "0010001001101100", 
	 "0010001001100000", 
	 "0010001001010100", 
	 "0010001001001000", 
	 "0010001000111100", 
	 "0010001000110000", 
	 "0010001000100100", 
	 "0010001000011000", 
	 "0010001000001011", 
	 "0010000111111111", 
	 "0010000111110011", 
	 "0010000111100111", 
	 "0010000111011011", 
	 "0010000111001111", 
	 "0010000111000011", 
	 "0010000110110111", 
	 "0010000110101010", 
	 "0010000110011110", 
	 "0010000110010010", 
	 "0010000110000110", 
	 "0010000101111010", 
	 "0010000101101110", 
	 "0010000101100010", 
	 "0010000101010110", 
	 "0010000101001001", 
	 "0010000100111101", 
	 "0010000100110001", 
	 "0010000100100101", 
	 "0010000100011001", 
	 "0010000100001101", 
	 "0010000100000001", 
	 "0010000011110100", 
	 "0010000011101000", 
	 "0010000011011100", 
	 "0010000011010000", 
	 "0010000011000100", 
	 "0010000010111000", 
	 "0010000010101100", 
	 "0010000010011111", 
	 "0010000010010011", 
	 "0010000010000111", 
	 "0010000001111011", 
	 "0010000001101111", 
	 "0010000001100011", 
	 "0010000001010111", 
	 "0010000001001010", 
	 "0010000000111110", 
	 "0010000000110010", 
	 "0010000000100110", 
	 "0010000000011010", 
	 "0010000000001110", 
	 "0010000000000001", 
	 "0001111111110101", 
	 "0001111111101001", 
	 "0001111111011101", 
	 "0001111111010001", 
	 "0001111111000101", 
	 "0001111110111000", 
	 "0001111110101100", 
	 "0001111110100000", 
	 "0001111110010100", 
	 "0001111110001000", 
	 "0001111101111011", 
	 "0001111101101111", 
	 "0001111101100011", 
	 "0001111101010111", 
	 "0001111101001011", 
	 "0001111100111111", 
	 "0001111100110010", 
	 "0001111100100110", 
	 "0001111100011010", 
	 "0001111100001110", 
	 "0001111100000010", 
	 "0001111011110101", 
	 "0001111011101001", 
	 "0001111011011101", 
	 "0001111011010001", 
	 "0001111011000101", 
	 "0001111010111000", 
	 "0001111010101100", 
	 "0001111010100000", 
	 "0001111010010100", 
	 "0001111010001000", 
	 "0001111001111011", 
	 "0001111001101111", 
	 "0001111001100011", 
	 "0001111001010111", 
	 "0001111001001011", 
	 "0001111000111110", 
	 "0001111000110010", 
	 "0001111000100110", 
	 "0001111000011010", 
	 "0001111000001110", 
	 "0001111000000001", 
	 "0001110111110101", 
	 "0001110111101001", 
	 "0001110111011101", 
	 "0001110111010000", 
	 "0001110111000100", 
	 "0001110110111000", 
	 "0001110110101100", 
	 "0001110110100000", 
	 "0001110110010011", 
	 "0001110110000111", 
	 "0001110101111011", 
	 "0001110101101111", 
	 "0001110101100010", 
	 "0001110101010110", 
	 "0001110101001010", 
	 "0001110100111110", 
	 "0001110100110001", 
	 "0001110100100101", 
	 "0001110100011001", 
	 "0001110100001101", 
	 "0001110100000001", 
	 "0001110011110100", 
	 "0001110011101000", 
	 "0001110011011100", 
	 "0001110011010000", 
	 "0001110011000011", 
	 "0001110010110111", 
	 "0001110010101011", 
	 "0001110010011111", 
	 "0001110010010010", 
	 "0001110010000110", 
	 "0001110001111010", 
	 "0001110001101110", 
	 "0001110001100001", 
	 "0001110001010101", 
	 "0001110001001001", 
	 "0001110000111101", 
	 "0001110000110000", 
	 "0001110000100100", 
	 "0001110000011000", 
	 "0001110000001100", 
	 "0001101111111111", 
	 "0001101111110011", 
	 "0001101111100111", 
	 "0001101111011010", 
	 "0001101111001110", 
	 "0001101111000010", 
	 "0001101110110110", 
	 "0001101110101001", 
	 "0001101110011101", 
	 "0001101110010001", 
	 "0001101110000101", 
	 "0001101101111000", 
	 "0001101101101100", 
	 "0001101101100000", 
	 "0001101101010011", 
	 "0001101101000111", 
	 "0001101100111011", 
	 "0001101100101111", 
	 "0001101100100010", 
	 "0001101100010110", 
	 "0001101100001010", 
	 "0001101011111110", 
	 "0001101011110001", 
	 "0001101011100101", 
	 "0001101011011001", 
	 "0001101011001100", 
	 "0001101011000000", 
	 "0001101010110100", 
	 "0001101010101000", 
	 "0001101010011011", 
	 "0001101010001111", 
	 "0001101010000011", 
	 "0001101001110110", 
	 "0001101001101010", 
	 "0001101001011110", 
	 "0001101001010001", 
	 "0001101001000101", 
	 "0001101000111001", 
	 "0001101000101101", 
	 "0001101000100000", 
	 "0001101000010100", 
	 "0001101000001000", 
	 "0001100111111011", 
	 "0001100111101111", 
	 "0001100111100011", 
	 "0001100111010110", 
	 "0001100111001010", 
	 "0001100110111110", 
	 "0001100110110001", 
	 "0001100110100101", 
	 "0001100110011001", 
	 "0001100110001101", 
	 "0001100110000000", 
	 "0001100101110100", 
	 "0001100101101000", 
	 "0001100101011011", 
	 "0001100101001111", 
	 "0001100101000011", 
	 "0001100100110110", 
	 "0001100100101010", 
	 "0001100100011110", 
	 "0001100100010001", 
	 "0001100100000101", 
	 "0001100011111001", 
	 "0001100011101100", 
	 "0001100011100000", 
	 "0001100011010100", 
	 "0001100011000111", 
	 "0001100010111011", 
	 "0001100010101111", 
	 "0001100010100010", 
	 "0001100010010110", 
	 "0001100010001010", 
	 "0001100001111101", 
	 "0001100001110001", 
	 "0001100001100101", 
	 "0001100001011000", 
	 "0001100001001100", 
	 "0001100001000000", 
	 "0001100000110011", 
	 "0001100000100111", 
	 "0001100000011011", 
	 "0001100000001110", 
	 "0001100000000010", 
	 "0001011111110110", 
	 "0001011111101001", 
	 "0001011111011101", 
	 "0001011111010001", 
	 "0001011111000100", 
	 "0001011110111000", 
	 "0001011110101100", 
	 "0001011110011111", 
	 "0001011110010011", 
	 "0001011110000111", 
	 "0001011101111010", 
	 "0001011101101110", 
	 "0001011101100001", 
	 "0001011101010101", 
	 "0001011101001001", 
	 "0001011100111100", 
	 "0001011100110000", 
	 "0001011100100100", 
	 "0001011100010111", 
	 "0001011100001011", 
	 "0001011011111111", 
	 "0001011011110010", 
	 "0001011011100110", 
	 "0001011011011010", 
	 "0001011011001101", 
	 "0001011011000001", 
	 "0001011010110100", 
	 "0001011010101000", 
	 "0001011010011100", 
	 "0001011010001111", 
	 "0001011010000011", 
	 "0001011001110111", 
	 "0001011001101010", 
	 "0001011001011110", 
	 "0001011001010001", 
	 "0001011001000101", 
	 "0001011000111001", 
	 "0001011000101100", 
	 "0001011000100000", 
	 "0001011000010100", 
	 "0001011000000111", 
	 "0001010111111011", 
	 "0001010111101110", 
	 "0001010111100010", 
	 "0001010111010110", 
	 "0001010111001001", 
	 "0001010110111101", 
	 "0001010110110001", 
	 "0001010110100100", 
	 "0001010110011000", 
	 "0001010110001011", 
	 "0001010101111111", 
	 "0001010101110011", 
	 "0001010101100110", 
	 "0001010101011010", 
	 "0001010101001101", 
	 "0001010101000001", 
	 "0001010100110101", 
	 "0001010100101000", 
	 "0001010100011100", 
	 "0001010100001111", 
	 "0001010100000011", 
	 "0001010011110111", 
	 "0001010011101010", 
	 "0001010011011110", 
	 "0001010011010001", 
	 "0001010011000101", 
	 "0001010010111001", 
	 "0001010010101100", 
	 "0001010010100000", 
	 "0001010010010011", 
	 "0001010010000111", 
	 "0001010001111011", 
	 "0001010001101110", 
	 "0001010001100010", 
	 "0001010001010101", 
	 "0001010001001001", 
	 "0001010000111101", 
	 "0001010000110000", 
	 "0001010000100100", 
	 "0001010000010111", 
	 "0001010000001011", 
	 "0001001111111111", 
	 "0001001111110010", 
	 "0001001111100110", 
	 "0001001111011001", 
	 "0001001111001101", 
	 "0001001111000001", 
	 "0001001110110100", 
	 "0001001110101000", 
	 "0001001110011011", 
	 "0001001110001111", 
	 "0001001110000010", 
	 "0001001101110110", 
	 "0001001101101010", 
	 "0001001101011101", 
	 "0001001101010001", 
	 "0001001101000100", 
	 "0001001100111000", 
	 "0001001100101011", 
	 "0001001100011111", 
	 "0001001100010011", 
	 "0001001100000110", 
	 "0001001011111010", 
	 "0001001011101101", 
	 "0001001011100001", 
	 "0001001011010100", 
	 "0001001011001000", 
	 "0001001010111100", 
	 "0001001010101111", 
	 "0001001010100011", 
	 "0001001010010110", 
	 "0001001010001010", 
	 "0001001001111101", 
	 "0001001001110001", 
	 "0001001001100101", 
	 "0001001001011000", 
	 "0001001001001100", 
	 "0001001000111111", 
	 "0001001000110011", 
	 "0001001000100110", 
	 "0001001000011010", 
	 "0001001000001110", 
	 "0001001000000001", 
	 "0001000111110101", 
	 "0001000111101000", 
	 "0001000111011100", 
	 "0001000111001111", 
	 "0001000111000011", 
	 "0001000110110110", 
	 "0001000110101010", 
	 "0001000110011110", 
	 "0001000110010001", 
	 "0001000110000101", 
	 "0001000101111000", 
	 "0001000101101100", 
	 "0001000101011111", 
	 "0001000101010011", 
	 "0001000101000110", 
	 "0001000100111010", 
	 "0001000100101101", 
	 "0001000100100001", 
	 "0001000100010101", 
	 "0001000100001000", 
	 "0001000011111100", 
	 "0001000011101111", 
	 "0001000011100011", 
	 "0001000011010110", 
	 "0001000011001010", 
	 "0001000010111101", 
	 "0001000010110001", 
	 "0001000010100100", 
	 "0001000010011000", 
	 "0001000010001100", 
	 "0001000001111111", 
	 "0001000001110011", 
	 "0001000001100110", 
	 "0001000001011010", 
	 "0001000001001101", 
	 "0001000001000001", 
	 "0001000000110100", 
	 "0001000000101000", 
	 "0001000000011011", 
	 "0001000000001111", 
	 "0001000000000010", 
	 "0000111111110110", 
	 "0000111111101010", 
	 "0000111111011101", 
	 "0000111111010001", 
	 "0000111111000100", 
	 "0000111110111000", 
	 "0000111110101011", 
	 "0000111110011111", 
	 "0000111110010010", 
	 "0000111110000110", 
	 "0000111101111001", 
	 "0000111101101101", 
	 "0000111101100000", 
	 "0000111101010100", 
	 "0000111101000111", 
	 "0000111100111011", 
	 "0000111100101110", 
	 "0000111100100010", 
	 "0000111100010101", 
	 "0000111100001001", 
	 "0000111011111100", 
	 "0000111011110000", 
	 "0000111011100100", 
	 "0000111011010111", 
	 "0000111011001011", 
	 "0000111010111110", 
	 "0000111010110010", 
	 "0000111010100101", 
	 "0000111010011001", 
	 "0000111010001100", 
	 "0000111010000000", 
	 "0000111001110011", 
	 "0000111001100111", 
	 "0000111001011010", 
	 "0000111001001110", 
	 "0000111001000001", 
	 "0000111000110101", 
	 "0000111000101000", 
	 "0000111000011100", 
	 "0000111000001111", 
	 "0000111000000011", 
	 "0000110111110110", 
	 "0000110111101010", 
	 "0000110111011101", 
	 "0000110111010001", 
	 "0000110111000100", 
	 "0000110110111000", 
	 "0000110110101011", 
	 "0000110110011111", 
	 "0000110110010010", 
	 "0000110110000110", 
	 "0000110101111001", 
	 "0000110101101101", 
	 "0000110101100000", 
	 "0000110101010100", 
	 "0000110101000111", 
	 "0000110100111011", 
	 "0000110100101110", 
	 "0000110100100010", 
	 "0000110100010101", 
	 "0000110100001001", 
	 "0000110011111100", 
	 "0000110011110000", 
	 "0000110011100011", 
	 "0000110011010111", 
	 "0000110011001010", 
	 "0000110010111110", 
	 "0000110010110001", 
	 "0000110010100101", 
	 "0000110010011000", 
	 "0000110010001100", 
	 "0000110001111111", 
	 "0000110001110011", 
	 "0000110001100110", 
	 "0000110001011010", 
	 "0000110001001101", 
	 "0000110001000001", 
	 "0000110000110100", 
	 "0000110000101000", 
	 "0000110000011011", 
	 "0000110000001111", 
	 "0000110000000010", 
	 "0000101111110110", 
	 "0000101111101001", 
	 "0000101111011101", 
	 "0000101111010000", 
	 "0000101111000100", 
	 "0000101110110111", 
	 "0000101110101011", 
	 "0000101110011110", 
	 "0000101110010010", 
	 "0000101110000101", 
	 "0000101101111001", 
	 "0000101101101100", 
	 "0000101101100000", 
	 "0000101101010011", 
	 "0000101101000111", 
	 "0000101100111010", 
	 "0000101100101101", 
	 "0000101100100001", 
	 "0000101100010100", 
	 "0000101100001000", 
	 "0000101011111011", 
	 "0000101011101111", 
	 "0000101011100010", 
	 "0000101011010110", 
	 "0000101011001001", 
	 "0000101010111101", 
	 "0000101010110000", 
	 "0000101010100100", 
	 "0000101010010111", 
	 "0000101010001011", 
	 "0000101001111110", 
	 "0000101001110010", 
	 "0000101001100101", 
	 "0000101001011001", 
	 "0000101001001100", 
	 "0000101001000000", 
	 "0000101000110011", 
	 "0000101000100111", 
	 "0000101000011010", 
	 "0000101000001101", 
	 "0000101000000001", 
	 "0000100111110100", 
	 "0000100111101000", 
	 "0000100111011011", 
	 "0000100111001111", 
	 "0000100111000010", 
	 "0000100110110110", 
	 "0000100110101001", 
	 "0000100110011101", 
	 "0000100110010000", 
	 "0000100110000100", 
	 "0000100101110111", 
	 "0000100101101011", 
	 "0000100101011110", 
	 "0000100101010001", 
	 "0000100101000101", 
	 "0000100100111000", 
	 "0000100100101100", 
	 "0000100100011111", 
	 "0000100100010011", 
	 "0000100100000110", 
	 "0000100011111010", 
	 "0000100011101101", 
	 "0000100011100001", 
	 "0000100011010100", 
	 "0000100011001000", 
	 "0000100010111011", 
	 "0000100010101111", 
	 "0000100010100010", 
	 "0000100010010101", 
	 "0000100010001001", 
	 "0000100001111100", 
	 "0000100001110000", 
	 "0000100001100011", 
	 "0000100001010111", 
	 "0000100001001010", 
	 "0000100000111110", 
	 "0000100000110001", 
	 "0000100000100101", 
	 "0000100000011000", 
	 "0000100000001100", 
	 "0000011111111111", 
	 "0000011111110010", 
	 "0000011111100110", 
	 "0000011111011001", 
	 "0000011111001101", 
	 "0000011111000000", 
	 "0000011110110100", 
	 "0000011110100111", 
	 "0000011110011011", 
	 "0000011110001110", 
	 "0000011110000010", 
	 "0000011101110101", 
	 "0000011101101000", 
	 "0000011101011100", 
	 "0000011101001111", 
	 "0000011101000011", 
	 "0000011100110110", 
	 "0000011100101010", 
	 "0000011100011101", 
	 "0000011100010001", 
	 "0000011100000100", 
	 "0000011011111000", 
	 "0000011011101011", 
	 "0000011011011110", 
	 "0000011011010010", 
	 "0000011011000101", 
	 "0000011010111001", 
	 "0000011010101100", 
	 "0000011010100000", 
	 "0000011010010011", 
	 "0000011010000111", 
	 "0000011001111010", 
	 "0000011001101110", 
	 "0000011001100001", 
	 "0000011001010100", 
	 "0000011001001000", 
	 "0000011000111011", 
	 "0000011000101111", 
	 "0000011000100010", 
	 "0000011000010110", 
	 "0000011000001001", 
	 "0000010111111101", 
	 "0000010111110000", 
	 "0000010111100011", 
	 "0000010111010111", 
	 "0000010111001010", 
	 "0000010110111110", 
	 "0000010110110001", 
	 "0000010110100101", 
	 "0000010110011000", 
	 "0000010110001100", 
	 "0000010101111111", 
	 "0000010101110010", 
	 "0000010101100110", 
	 "0000010101011001", 
	 "0000010101001101", 
	 "0000010101000000", 
	 "0000010100110100", 
	 "0000010100100111", 
	 "0000010100011011", 
	 "0000010100001110", 
	 "0000010100000001", 
	 "0000010011110101", 
	 "0000010011101000", 
	 "0000010011011100", 
	 "0000010011001111", 
	 "0000010011000011", 
	 "0000010010110110", 
	 "0000010010101010", 
	 "0000010010011101", 
	 "0000010010010000", 
	 "0000010010000100", 
	 "0000010001110111", 
	 "0000010001101011", 
	 "0000010001011110", 
	 "0000010001010010", 
	 "0000010001000101", 
	 "0000010000111001", 
	 "0000010000101100", 
	 "0000010000011111", 
	 "0000010000010011", 
	 "0000010000000110", 
	 "0000001111111010", 
	 "0000001111101101", 
	 "0000001111100001", 
	 "0000001111010100", 
	 "0000001111000111", 
	 "0000001110111011", 
	 "0000001110101110", 
	 "0000001110100010", 
	 "0000001110010101", 
	 "0000001110001001", 
	 "0000001101111100", 
	 "0000001101110000", 
	 "0000001101100011", 
	 "0000001101010110", 
	 "0000001101001010", 
	 "0000001100111101", 
	 "0000001100110001", 
	 "0000001100100100", 
	 "0000001100011000", 
	 "0000001100001011", 
	 "0000001011111110", 
	 "0000001011110010", 
	 "0000001011100101", 
	 "0000001011011001", 
	 "0000001011001100", 
	 "0000001011000000", 
	 "0000001010110011", 
	 "0000001010100111", 
	 "0000001010011010", 
	 "0000001010001101", 
	 "0000001010000001", 
	 "0000001001110100", 
	 "0000001001101000", 
	 "0000001001011011", 
	 "0000001001001111", 
	 "0000001001000010", 
	 "0000001000110101", 
	 "0000001000101001", 
	 "0000001000011100", 
	 "0000001000010000", 
	 "0000001000000011", 
	 "0000000111110111", 
	 "0000000111101010", 
	 "0000000111011110", 
	 "0000000111010001", 
	 "0000000111000100", 
	 "0000000110111000", 
	 "0000000110101011", 
	 "0000000110011111", 
	 "0000000110010010", 
	 "0000000110000110", 
	 "0000000101111001", 
	 "0000000101101100", 
	 "0000000101100000", 
	 "0000000101010011", 
	 "0000000101000111", 
	 "0000000100111010", 
	 "0000000100101110", 
	 "0000000100100001", 
	 "0000000100010100", 
	 "0000000100001000", 
	 "0000000011111011", 
	 "0000000011101111", 
	 "0000000011100010", 
	 "0000000011010110", 
	 "0000000011001001", 
	 "0000000010111100", 
	 "0000000010110000", 
	 "0000000010100011", 
	 "0000000010010111", 
	 "0000000010001010", 
	 "0000000001111110", 
	 "0000000001110001", 
	 "0000000001100101", 
	 "0000000001011000", 
	 "0000000001001011", 
	 "0000000000111111", 
	 "0000000000110010", 
	 "0000000000100110", 
	 "0000000000011001", 
	 "0000000000001101"); 
 

end DDS_constants_pkg; 
