

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
g1WA8VSKrKaR8FNxaZhO7xwQ1AuSq2XfGW/Qob1EGM1eOp/C7nueVpgo94v8J5uGPaQKqd6kfYya
m+/Y3uxo+w==


`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Pu2n0nCiuVDDFE8CzoDoOjwZp/WID/e6m6DQC3SyqRSsbuwi46xXY16nPXUjhw5kf+V1TwmkBF9i
yG37oRNjwmJvXpDuTO0XV7sp+XSRqDaGUe2pRkpRBVBU9P3VV/IST113kZ3am41lRlJljYp63lHV
Vdqryd6Kvm7Nnmls7W0=


`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AWYIBGoZpXrmXMqZZuDG8Z9rmprtBozCVQ3s5hRfiCNveIF7IQfYW3QcouzsExTjEljAUOYqSWIA
ZxjaxjtqmIXnozCa3TDXnYopjqBNNh98OjjEm+aKt0KQUGl7TboeJFNIuOZTBvg4XkBnu1olCazS
vlVdsOKMgzdkUo+rqq6YWwLZOD9mWVk0KTVF33wZHYV+5YlKhwkF8dHO67W89Li8er38ELkHVclN
7Xs+cDR4EX93OBOrQmANjgH0ggrROY3MJITcehCOK83VaeySfrKLrqKlcWpXqdp6T6vibEe3et1O
pG+et5MtIWoEi1yt+W3qZS344mwAh52+ybVasQ==


`pragma protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
g6bvjSvJ33u8knsw3IZCHpiZrDz4KX7MzVtz3VpD/Fq0RYDpUvUcUFPvoiPL3jExQSuEUc0Aq2yg
xmubv5Pv+b6uycpQSt3GN8QtFfv3xA0xM09bctvjmD/J70V1ZwTFfUhFn/KnXwKt0MgiLAT3uy34
1u4/ZSEUTSxO0MCysMBwQhiobY6DBOQ3mHD3wAw4lFosW6S+AhrUNmSBv1EPxN0N2WY3nF3eTibF
neBQshuXKow5C16okE/MLogv5yqYEo6aV7E6aQGWon2Hl7KRVLHVcfiqn/Z8l2VaVSPxylmdvLCV
SB1keK9AGFPpb3uMR172fw1vZm88a5NJB4XO5g==


`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
GSC8Q4Y0okKWGHWMU4J51XV+Fp0ojryrkqw8EEkQFsdx/xfWuXFtV37ndIDMp/i+0GAIIFK+m6BC
fkdQHMVu2bss7g0J3nO37fGZRLPKrdlXghl1AjlQy+Y/TiuroOwyvs030a7B+U3A70WGnFe+/w1D
hISURUJkh2gQi2aOCsuKW1c3+k26rSmn5QruazNrIHmGG5jwEKsPdgsEdkTI4n5kPRVocW4kiLGs
mQh2/QI0LQd9Tydq8rBc8DmOFjB1VHyUZO3CdbU797YR8Edx9/o+qy3cej2bw6rYOnHiWe6XhTur
aL6LvYo5Nc0misaf1+6LL+bnZi+vng6ec5fq5w==


`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
cLTTkVlQulW7iOySvGIvfdifPC5X3pSfOgLcUFhU78V6Tehu6ogGn4KXzHllDPp6IRLgb1oZNQmP
WHSVVLgJQF+gI9RHoda864s4uG8VdB0stSlgQz0NIlfvci++wBDa+4+EG0g7svbVj2R77DrxZvqC
24ua9OVOM7I/1Oi+PFE=


`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
M+WFZmxctI4CpxmlgnXJJWnslwOutoAvtZu5bdnqi3mO+DxDLgDDGpn59ids7G1G/FhgnDA54WpO
FLuJ5lluv5iaXjtZKvvdLGFq89MOmL1+ePrHT80dyoWq2yUvQfi2QQSdyZImABhQnB5kCyCSlg65
06f66h0aASv7ooP+XrxLR90ziTXJGeAJ+da29nymGLuandzJARo3KEpPqi5IwbBRHCsvxlsU8Vdg
V2aOPLvkZIUY5PZ+ZtVmQPnNDUie5F/umbLRumB1hid51Pwr/RHxdIHM8WDQgO/9HAYbZrI7O0Wj
FSY8Afp7d2yVPf11pzYQDEm15lWUbCdQC4WOtw==


`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 220608)
`pragma protect data_block
svFl2EBzXWKFBsDYBMcKma43DgPjpum/OhdssnGStTFJU2/iSxRBu9ha6BegWPMISJTKJEI4yK1K
1etuDgvNPqkzT5GI+giPEcbEPD/kM8XOIVr3inOJO1dg1KOyUVQkqeMkUjYxhn1bAyg+PGycqD74
9yMAy+DxXDPnQSryMyB1z3WPXM8VGMk4qYT7UIEmGwaxcF1Os5Ybkoc5G1d3BZbfviFZiUTqCxch
EuGbnFDH9mq5Zxqe0+oZf72X4Bfhxwk/ZB+XaE3d6BFyB5iiux5Jx1kcQ3Ha2k54MSnIgs6hNv6N
/eD8eDuVESGKEPxeBVHXNnErnKExDrjH72QZLWXDwgvO8D3SYkSHiy9/76rej5zi/wFVKCrg2hSX
cMAbpd2wk1cLjxgOWUdoOIXoKXqEjO9Gm+o6VcC9Xmq/aa23x2K6SxutMCys5c5rwQP9N+60OhH1
CQHxpswN/1y12ud/gxSvAYVcTMZC58hnPlfLW2ABfkmuO03xs3WYwLjg/uLZ1IK8zoTddUWYJtCk
16HolRDT4gej3d/SneFCwBDKNq+r+r9KFjW2xFu1hsHfhvTjI19AMQIr/zGM5cKi8LMUiEkKIM9l
6OOY8tqm21IrIPXo463jcIqvqCIN8br3dEZfeN/B4I/5oU39qM0UvceEmcqtJIVLH50rOhCmOJQc
ZQKKS7uemLH75o3MN4EFTcjyxxKq/sHv/5HV5oTx3sZlKkVgk++WnJeKrzoHHwceRSyRXWm1aBUy
lSjOXKOj7i8q2h9d4l53fVtssHZQBvOVfz+Q8V11RjPyCKbUVF7Hc03H7EHFmijL6UwVDfSSfe99
CHkqDTQsK3/c7lknYmHiBZOL10kgz2uu6A75oYL84yGoOySgel6vk3eBTWQr7q25tjgbIF6QTxPd
4UK029WxhfYFdj/Avq8vkZhlt6iGL+eywPeDO0KootBVLEhEDPznr7CQ5f4XFcGqxRTskaXehMTE
Sjxb+LTTIZ3obmfZDniG0iypdOfSnZoGHQFHr5zg0RHqzhST8e3ecb9xP5KAvo5JzPmQRZ4fgtQn
v6pksXuulpunIy+Bd7h+wBoUSd1Z1dS6zOr1bCWj/z12UwKdu5lTSI5Pzoi+3OBIxf7P0mVJnpa2
9iwKdTNYvkNZNYPHmUr9HvxC1H1R/y1OuoqbKT/KgBIH35B3cnCbSYo/gGY7ADGy4ZcWiEUny9MG
AU7THYNXGm9Z/zVpz5q632uQenPIm9lgJXnvzG0nKq/d7xFmi9+lyT1FmAM9mWdlryfA3jh+QjQQ
0dGZtZ5k9NchniLIQl3GqKamUHC3WvP061h1vMfEt85nIwVw88wy+iPYJZeSuFkZm+3Qh1PnaSBM
kJFLM7zBg7n9b7m8zFZhqXBCPXtOA1ggk3BPDGTpKWDwlVQAr2l/8lwGtwLTmphQKRZrtUvGjYEW
FJUQOOmpaB+WJXIKtYGVYZcfUQQfPPSLJZvKkAizN5WH9+8n2+vA/a6YFxrn6N7boYh4Kw0DhIg/
aC0zEhe2Owidvf75YzVCPq6R+JF1J7PxpvpWxisIYxFWwpk8BPDInqSh8qXOP9jnURjhgZVINNRF
E0oNjnSg5+RmfXQV/U4UruhJU8KfHTqxGSyV3hMc6ea0ajXHUf2FuJtKLuvG9em3aDIpK/UcbgtF
fAZFNXNQJ8NVHpaWs23Z0k+PUgOgjVsNpVT02yS3vMPUsdZ9jGEfQM2+F6g9WdZarKH8zBTZnVA8
w9I/0jLhcdULdQaVzyYgDDDfHnnCwFVbWXbz70Wqs4Gjbfr9eG5JsA6pgOMM+HMFxHnw30kFi9go
cCLgY5ReshYOUY6576BZVhbe1uXCmSxr+8yvKayFtG30n8I/m3nze/dthHBnSpL85fRgd5eWsfpH
UrxvRrUgZ6h4UZK0mmQBnlnKrbroCsWilukQi83xIB4tgSbm5c2vETPW5vaZB7TGO0PAUap7TNXm
++RLhsgneybbu7AjW6SMjfw9VCJzpSxqG1AF40uwmteZZmGNV+DT7Ey1KZ6sAHZJmFEcjMytMoh1
BMZXcoR/1GDDNjLUEVOi9BFUE/XGyyw0FKYFi4wbVqO/1mRFatDG88rxFQyrqR5G83hlUksIettj
XJppEX+QsnbPOx0SEuDRjLhWwlIIr7ahPFtZktrW0MEXCZhix0x1PYl5B896MIoQoDzKXINZ/6Vj
VEiF92PnkDV8E0r27mlo+O023fOZzpAlIIT3lvTbk1bnRdtAWf0iLmFBPyRxZ3Z14ckoY5/Mnl76
bYZnkkC+mkR38hUh4KOfly2XXgeZQ+5Pun9+ybLt4251ODzjKB5WLzLVSxn06JL+De1Mt7bUw5r4
Woj52gN3sRB3jcLFOFFxCe61UL0IrrIiHnzUz6lbT5icxmIkZpodLkTDIGhohI/MiRPsazBz+ZU4
qvMuzAkVGZzO4aogwirV3tTu4issmHUDO8Y8JS8RduKfnJydlsjd5SN/VVZ+H18gEUytaD1xETHT
tl2rQRrNA7K4Q/I0yLB4O8UDftc90f6LzT0tauw1pHiTPQda0T3ioBvGRi71oD6ttKNKnjgrSVhb
QxAsYusdR156hu2Y56xjMJpcSWaGTanvp4BJ081XJCupw0j1AmsuR16ZUzyjwt0yRLSIsYdCoMzY
WJufT5xbJ2hgqNj99DlHtONFwjahN0zytDy5GwinL1lEQ8dAUkCbChAjI44vef3iZZVUKtCl3UCI
pGBkbPh5KHkLPixXwPFKTBBV/VxinePC9vuOIzJgutbDWloxL4/qFyY6NLTvBIFhwjuS4ozDzmQO
RLAQNIadASnX+aLK1YBi9fU4ltW9sD1bQv5aghUPaFD5m0Xl/S0eBS/eB/rnsCwTxMPg3lhJ+20h
gSWnkCKIdWMdQPiCyYPGXOA12iDbt5Cm4L34H6qmVdeHLj5QqGOpMh4sTMmiyks6OLspa/A+ck2j
jOn445z4KoFGaaST0w/yq7ZgJP1OtgwhW25eeeAlAZCXw5lHfgHm6XuenDWemYgOTyNuGEYkAPeR
B8e4JbX5mNPRsLiEDeg3qsqydKIQDW2B+GRWwV4CWWjtPwzVTY+O97yR1iS0xSq871EoLuiBwkvU
cZCFOj0vEksyAo8ypeRhfI2ZVEkhhs0fYT21kkHgX7LCakPREtkKIKSsLmCAVb6Dvm3KudteYdWp
fPUX2a4KRmUai296v+g7i2g+jgDhx0ui5LpVtvHT7IIshJ9tiOqdAyDeFHHP18GeVjB5I64iRWWZ
0dMOKKJfRqQ0WeETWt+9s7ZHtQdoQ0Y9+6DLjxJXm1pT56OovmpPK0GKwg4+ow4GkeEOIDCHHPo+
JBBg+/Dlq3nJ3hoy0ikMxYx0PL7mP4d8dG74P5fkWMpc0yEAmuMm5iEwi5lOLLXGONjIKLRbUwHw
P3ZACosA0pkrphS09GnDnkdOU3gCkX/aBt+S7z6C102yAcyCQoc2VVwoMHDnQIfo7Qaa+NkR1Vrx
2a/bCEFKqVQR/5rzpsDXT4qOAjfpaNemDUJ50vDm8AunK3TDMTir1zZQegRGYwjhTps2zyALhjZZ
n3NxP3WQrI0+yHBIPOcfkPeFDJtSl7C/I+/2ebYmrQAwWEZmWQF2QWGkdpE5d4KyztU2acQ+7SCo
5PzVBw3Zaok/s3xU9L8A/Wmu5kuZfwPbbCjiL1a6AxE6ATeR2YIJtBC3kK8UUJtTRiaHPLe8M1K3
jjrnI/b7UiSEgvWZJiXwAh9MeGXVQasyW+vPRcQzOsboud+XjiiKuRQR4blDGq1p/DQZ9IUbydOy
p0sp+rr58a8lmWmvlUTtqKAVA0DFirJIPfh1fKJp8TizVTfW+M2uLDXcTzs8PNN8Zx8OgondV5q8
bNK0h8BcrVtHvoDBBUgIUcnfV5cglw0seL3u1BJ4hSKYoi1D5z0AqMrAQATrynBe6banMrCIIOZh
huq1yjOVK3xrBQY4vXvS7IDgUxkgN9PmnDMov1jDWppd0jbcWOIUHelTlS/MKAvJ5/KVq5RUcKsT
bUgs/tbTpD2CpQRcPnTENS4MNLkc+qJSaHJ32FCmMdJLqO/Sv6hQBSrQ41bu+O2ELKGEJqN3R4B/
ER54O9qdw454X1Os6as2gqtvNAUfYZ+0vLxWaoWuA4ByK991g0RO0Al1GHUE80pBE+YKW4P4NecE
fOXagYcDWAD6L9Y622N2TWldc7cqirVYl9+qRQdLOFEdA1m+b0kOTDbSLrCh92x/+2PKk6ltKJov
YVoZB9FZG0IiVVT9xpAZOFlRtMwUA1vI815ITqLvNdOaEyApFAMZYVGGIYqNggRF9Cfo32KlCofP
dmF2fFkzkJuFJ/7e60B9JD3ADIMaGRvfqEa6miSgqBfYXNh7cR7+VHiAgA4KJ5hvFNTN2S8lk+Il
4qkdyfU3xERpmJW+flB4zKwZlquCzly+IbzrevSkCI2K6wqqFiqByPQ1+/iWnWHDbHKs5U0/wWCO
yKi/DcePNXGF1d3ANtT6w8hzU4HMgjcD/Cjfx6xlq5WH1mUf6xt2JmXCVK0bYbtL/t/fH3lQc24b
98qfaNFvgTJXZhH9kuzXFC7NhJ4462OQarVeuMj8o7ea2BZBAv5NFlyaJH1rGBfCffjRcFC6Uzqj
KJv1SRjA7GOEQtR8dQPDwFmA9uGCGmWlQuc03dqdFJvUVJh5NwcUpvRik8e9EJiEFEFzK0T6WWB7
lsvMPR/bxHwlI33Wt58bh8HpSdHO7SwcucEsbTtsjwmmgbNDcEay7MdH6fCRpGhiA+YgW5XLTur9
t/HhUkyS+eAx5/vI1lmnjtUCT0Scu1/NQHXQa0Vz0fIBjk8D8/kcoayfxH6ZLi34UsE9SEI/c3wW
4go9rX3AU2lTkm5I2mu6ymhKT9D/W+jr34lIQgtNrVdDokkHAAVzgHcon52kO5cZrVvqMrKpn3uj
pwj4RnI58pnXLQhrphtOP4pepemwqypqDlVkksNsQ5wTnDGkYW/K/TDW1HKwZG9dNqeVxha+tBjX
EIpCvibc1C+6UbUcOo6rRKYY/kUUb233EDly6i6z6Fwi7TqXOX32GT/5SPQuQAXh1nHPyIkGh3EJ
HXyUJ/iM/hLYU5bVZCfZp3YkNOuAYbe4gN4C2szaiQuRucbZbe3VBAxNJwlle68qn+nPpJQbOdc6
/2Q1O7vUD1SmohjbbeD/Ubm/4qVDsoSZOSuF8hETH89Wa+IYXRvIQFAPyzRFEndHCNtrJCD87sHG
84D9myzzJCwuN2iLnK0maAQeD+uBqngWq57k7/T//xkzK7aPENZbiwNTZ9k9mW6zwi3lG+cpCdMG
2RTpKqT+AliJc33/9QIEO5CIFy83N65vyyVuG/ycnLH+KrWeWK3Os7OV05PjKGUDPhReW/BYiwEv
tT80kTNa02VTZ4TA4HpCtGgJBwMgOrIh12GZARaPLcGzGecL/WqOyTLOTU873fTBw6SIN2cyWmbC
7nyncW1nPv+kv+7yW0FFDQQPmL5E5PJo7XJ57QwM7SnGc1WT4gHm154BoZusZ9TUWdWbkEyPGWdC
WWpoSZmvnSppSuvnvwDkdg9pcz5aamSD1vP7MeU6mA2hvLD05930/Xm/eqZ3RAXg8cj9ERhov4gU
ompqxnm3eUyF0y9XvtrpFpjM3/thcODIqsagogYrVdo1JZcA1Vb3Xq98hO2+hNnk0xpQ1LLhasB5
MWqXNhBpbAD1RYPTq31o9qFnqAlOvQxSoG60fbMn3uq6pYIyMd5Edwts9CKnmftrX+okAvQpGnxz
/npdj65veMeMiNJyaPnjsmC2kmm/legh5wFHlrobIoDOM+KYe3jqpZbPkOOOdWOwfVrqbXinor37
5ZBTTVjLl+c96Di0/ogHJLPAlR4F3a4zW3b4lT5Y+cNQUQ8nzEPaPXMtpDSN6ydUwOaOyxhqRhNo
EsKozGUW0HITXnk6tI3kRz1zU2SZsGsPT3rZ+3/qHwZf6jR4pwyGexfhQXFAhYVMdmfmAupP790j
ObBYpqaOytVMwddlGLWr9SI2mygV9nLBcPvjqbqH1AO+pXyPmmfIgurhdwUcKkRDkdfQVdXsSHHR
RtKXPDtBUG1TwSXuRUGK0lHD1JvVVq9gTsMVld2kUUDw+9mrOH/OP/m35FvRJevjFGC042UZEJXy
LSI1iI1Ri9aIFdyOkY7A00AI46NhO3p0JjU975U/3jJ/LLbuAkrFXQGncFYxXimS9typP15VF8Lm
AFC4IPuqO+PXdprMcnBQyK2SxBRv/Ve8UHuLVPZvHC5wlbwLnjKTPIWFkCIYY7zfhLax4YsXHLcR
b8rGIcbYzMwqHT8u5/pvuAhvhn1ZVlgrLEMJQUSGxFthEq2wcviqsbhWKhhuPheJ0Y0SN8UmROvL
rVbPfVpbVTG6vmBTK90RnEJgxCppSRonAm+2Tpgn4MM6dWdmyL3bbYPF3hFAkYUDP9sa6DlnZNZs
ASTx3x4Of3wrFIAUqiKhZOPDUgToyugB8qSFef6zzVHjlyfOVQXyri2kzmD3YMj4GTKZsPM8f/Yk
6hNDg1RDNqZwHfMbQzCDBsHHWCKdOJrp1hn9oXEJV3H40ovVuHsojZChW/yqkdFr05pb9AEDMJHN
k69tKoVwHS3W97bQ0RezOts4Ytr2yj02rtWAaJXf0dyoJLRJRzqWD500gdR+tEf8LOo8tgK68mM6
HsAoxlSNZLu+kN2h82nfEl71kr+O43OyIEv39LLwnKTAszFRICzAE7rqmU6z2Mp5OaOWA/ronowX
arKqa5Cta/jHdnXF7zO6RP6rEj/wfHoFSvouu3179Vu+havIIEPNsRe4QwVJ/0h7qi9MNBErxrUS
/1oNO5Smco/V2hqm2ZKUIy+H4qh8pjv8Qwn0xMnkhGDDKaeHSg65ujN2PNKeJmenQTFMwUnIo1fE
pYRMP9gNv3yNvIt+508zH3SBi041Xwc0UytoztVfP6bpahXbzWjMgEapIdkTYxCZbbm45QoaOpQo
xgwGk69YmnSgV/N2aKRzHRWGGlp68nhHaZk/4GHI2s0648loHVz8fhqXgG+jE6ybdD24F4tKczOr
IZuGwvP7v/CfBYzou2Rh9Cp0r81OIC/KNUHWSW6dU38J6F/3y0zaOMwRZzhl1+rZlDjeRd/Df01k
CBcHN3+TnVCAdJP2VQU9HJaZoZ3EZt6jvJVa3ZxDHKy30xhHbXmQREovv3cToaQSDg85gk70RXJh
pDnRUdL/xyrrUOTlgC9TGYQ12+lzQ4EWxueM7XmaJCEWIJNBNsl97nAnhkj5ys4Z3IFxMbqt881o
wpx3I6uNXSVVKjMITFsIlABASDVMgN0ylDuDjaj0pwy0UzlNMnrW3EYHNk0sPn7KdWOqCrHyKNwU
6Y3ZdteLsbTq8yL12iq8weAiMuz6571Fv9EwMlRa+/nc6EgFpVO0XMfVldc7Izwi2gteGis6N8c4
9nlRLfH9TlSs4eWancMP0I9c3T4pVP+AB8Tdr6D+vY3iUJxDrPOuqDj+ScsMq3BZw6lRCufDOZBR
hsnFNFGiMD6scM+jkirwy6zkjeZ3InvTednz/C5C9ld5dFc67OYAdgyZFDjihRrrSPSUv/4k+ANd
wRzbIHVYEq5JCRuJbCjpQrup5nq7bG0Hy79XigZ8VtNsKABp3AkQRLfGbD5Xss2Xts07R7VBNd8F
vykxmU0anjHEQMqpB6pe9ND4Tjx3VXM75Auwm8ySixL6ppT4ZTIoCUtBIaOc0eD9VhM8v4lmk1fU
DB04ynK4M8lm2mDIPFv3dUzbnq7StAwA6bWx1ZDomndpWaLt7ELp0G835G83wXr2AfHsSvDTNSwt
3uQyJNZ1WUa0ZsfRgdPfQchFJWKXqGprxFfnm9NaRF0C0TjMDc92+z1OdTaOijfvqY2eluTiQ8zy
lpalNbGwJrpur7/Y1fIac7ADUoQsPAWzse/FXff5AWlFSVvoifSEk9vjI9BBNxUNrUieZlSzSmji
w9uqm+yNPQ/thq20WSAnxVPjYXJM3nZ9qjWuI888O7/G/J7Q1DmtB9OSvF+IYMOz6ycL6wg/pXjc
xyIbcSbE53NS1GJl6C2Dzi58K8q2m2K0xh/M+SEMsmXZxuYJ6asBEnPb+5lATQM8YG56xtnziYeD
GOyN67qiKaJv+iH5pzQpE35mYtcUBL7HCKgH5aWqwuFe8PNKoClPR7i8jrzbBGADgKhNObw8m1kl
st1y/GmuRNDSAzOY8GFbiUHdeA0JW5uzEDVkzJjiqr3mTB+iVawS0udh5lA9lVzscdtbnkiU1IfH
YNffcsQCUwYIwkS9CJ3ydlASs6LuRO1LFLatZLUMzfPqo6pNVrpnCMUH2zP3YycfMQu9M1H1tIB9
DEjmyO9glhp6ig5wnpG8WW0UE87SffCWuFyOzPZZJFtV6yqRda5bpsppYPORhNDY+XHJHoBuwSSI
yUcrpVlg2eunmnUd4620k49Pmx5B8vXnJbLpDs8AKNQREcMC1YPg9dg1Sx2U9ya5flYhI6p750+l
/zegYYr2vQTUrFBYkPSxs0iLHFMyT26mk7599PrcFQzME1bQG68gUV5KGnRdw3OwYnzpS/t15wZA
tTYN/laTEilPGgON3QSVEhBsW577d+xqvXlNoQAlVy9JMJa8SPx1/AR7S11QafmyAdaxCKNEY+/4
wLAL+s4niZS6+6Czg7cSqIesjXzcYadTsQ4ODXxIQizX+KbsBYzaGH/Bae408clK2YdZUkvgBPGL
hsrP7DMeiRMkgllv74YGjI+vgxHQnf0uRNYx9G3QfyB1nDMiQr2ZF2xYpE9R/f7URQBb3SBfCY97
tRlQTTLHDMxjS6sITCtp3eaMTUwX+gdiZL2CZgnzgNnk97TtGSA9r54W5zK5YSeGTJdrt5UvexS3
w15EjVUIICWpk+vvPRk6x1xCdV+qjFZKKdSJSdcf220yqU6LZv+I/efHREqnRobODCdMZPXN9+ak
GwjIExiG0tZ5+KbwQloJ6ixoM4nJqM53G7wa24fKRdiW/wDe/bjZGq5nHSFhO1AHG90WFGoNWInL
3lH+bipLw/wFhvXdWr49TOawH5izV7bhH/UxIdyFm9OZE1/tS4wBh+Ik0MaYInD3ckOiwCB3tVbN
U3mG7VQgrGJETwrOc36K+v3s5eKwl74ZjJ1KWurbXD1sveCHbiiGFNaAL9SNn3XMHH49nQ3IHf46
tKJioRal4T8l1bz2301eTjzIKOoXNPdFKcbczY/hs9Zqn1o7DL5s+EgGE2BLu5JCX43wAlNyGDlL
x5Q1C7cIumThAFn8/BU9itbdcmNTxPNc+JbqzXBevcR9xg74dVUsksfQILaijVwa0Y5kRIJHv9hw
b/C5tTmcmeWPIAQ/toh/1WyC3m7/BlaGhimsxWFV0nBclkqK4tTXQpDGK/weSB9fJDd+Pztlr4u/
xzpfJYE3lcjHnTXwdZkk7Nm11WjP9CR6R2cCuKHaralmWvhE8EHx5zTsFpB2hMXw6KJJY5sRquL9
OyVnYonyPc6y3gWc5xeA1fQNXmfbq/g33qGetMIY9XnTITAtHvEvJUWsOp+8XBHfXLkzfIlhoZot
mTpjdsBlomwdcv2/PVARqNY/M6ej/fbwiN2JcMReuIkly72MF1Ny35Fe7GjebksXcBsbXqrMJtJA
Dys31oH0+lEjHevlaB2pl9iRnBq+0wt2cNTnK6/rUZ6bedamLUu9ccPpnrDtfH2gEoX7MnkNHyk6
pKJv/X0IGE9D3Auxp6rYBUGQx8wQnC/JXcOhVmDR2V46gM6+EKlFZHPh1jrhcjLQTfp56jKRgcyp
4310DTaRSxMjqIMkX2YiGKF1EUp+bpyW1pI4vgcIOfJDqCc/ZCJRFBSuUGvVKxCFWxgMW9WM/z+i
ItiKSAauGlFh+iL4AlSrt7ywRUdb7nUx5MFXq+ULaq+4CmdDvqpND9a9TzFjMopscbFIEa8P69e2
ETmzl2F323LgUBNii+pQ82HJ9p8jGC0fLZnzqCZhFd0x2TJEmjUCeLwjc2xjtMDYJy6WbZWD09ck
jlcC8WZrcHoE5pA8eHppMxjGTFS1XsYr97o+Rl4hiucTo7tC4IKGqbKg7EbY0XStJLum+TEtt2Ud
N8nhwDhzMFebk5dz/Eyjqp6jRbnoRK0W9cIHcqKBlMKFvrWlwqXvpsNKYZRRKOQmlEfEN57Yt0po
2WHf4O5Drv6N9IdCq9hxoXiNT1ii5RkIvvgJsYYqEwteR7c4kQC9fuOp5fx68YrisGEgOoxJfIw6
JRCveK6Ne/jxv9KhHCcbJamQaR0vs4AezYy6s6L+mWGwv4YHPh66hhzrJd5w8VA47KjTGSl0ZjAj
VQ54pSg+H4arsMcCiW+X7QOf23bXy7xIW5H44Helv2K6lKGVAIlWzjBI0/60YVBD2ZijccNw/nWF
Ou4++JhQrAHujByL0SXK2SwC5euD396b3NTpCEEq0SvMpCB8arD0uCGaCiRS2edLza0Co/Gw36AD
NRYmfHNiw5kA75bxM5AqgyZnkk/801zjIVdebIP8oCLNL7FIwXhaadx86qKUGua3KaazvhIgQYi7
15yFlVDpFsnvH9fvGNcGG0E0eYX3/0bjrWNy4AVctt5Sopk/dLOPKgKCYYQbPUI1eQht8/GSHJqy
c4dBJDuo0IVAHTt1QGUL04sHb3pB5ws9zQrcFtjtNAC+fZgSDVFHrjKePpVZn7Q4Nuw4vjRxVJax
8ZbXWGaYmsRk+StvOyT7See826xYy7BoHUFq9pQ8/j7tbROHtQBfxsno9sFHJAhQy0WSXhzFbKg5
SAnTaEqP4xBzyJIFAfEvPMEYoOPi+rtJavVeQzWqOGVOS/uDz8cjSnxB9SgPw6c7zIDO7ayEgs14
b7ngd6W4kqvIat5voh6m9uMFaeWBVhTUSUk4lqc/mlqNK+YV+NjyEMAdFEJJ5YDrtyd/h3DUhStt
IFU3GboQADPgBGxK0LmjI5sTbiRiyAZYiXYxj3yuZU2QLgcYNSVX5mCQf3nv7Czg1PTBs15o6823
+gn5krMD7bCVSZcsse7ZhX1WhgZtfZvZqTkjS7FbUdfVSBmoNfBotpYWKBiTsVOsOjP/j7gVyoy1
soXWLxYtR4dessRxz0JYDU6pH3uRyqNxxAJOc5LNVM2iJU4LYlYrZbdqCRsKhh/Xb29IKMxe7AUN
lxRWJt1pIJjRmr+EXFWbSldUdP4OQr41403wY3847eTkTyHMoLKdOZ+P4XeEmLTcGSdNWhL34ajw
5vfzqEGGMch44BksKXME3uyYn4Zug3cXrrlK3QxnAgaSLibYLTnEBh0ggePaLEy+h9yWbgYy/3Wy
7mVDYRz1xfHt0mQON1PSZsxUb6h1SCcoDxNIpIVuj0Q45AjJueM4nn4yc9zh7uAkxTs5IGwy+9Rp
0O3NIoQy5xZxk7plmJpFwsOkjVWvsqMpuU9mXciGHPC7BSFKbkvHdaQn5F0vNikA9Af1z5bDbZfc
MgvnTBcnyaj3cKui0Pp2Ggt7LoOSJXAI+I2XjqiqMLWHUTSX7Um/ivubDjQn1fm4hXzCuSgbHSKX
drdCT9f4tkuvY5NTDMQc0WjX/53ftEA1RqpLKBUGC6DaniG2UCLO1BqMFLMX8zWgBilyC/fb1jp0
qKD8Gtw90f9W8oMICL3oMVp7uGwHhHCtSzdNJx2+UxYquajFPuDNcrnPCf+eBQAS2ETgHAUwPHCD
/xqwIDhCkicG9ZGBJqmSHrzB+HIrqmi7x77A4Th5niKC1088B5NqRzavuV/TSuPOZelAZXPbMfwE
64EXdoaRLEsju9JxQFbJL2bAjPcmgC0sjAt1bqSP1T7W3OQeiaAZumtJYM7eP/5x/MkG9ddX9C+o
XfaHLp7vOfwhb6i3bS1u7ggLYMiLpa4TaepgAofsYeCSyWvpcjoPOOJMNiDrqKZDpZci/rEISAqR
9WDQou8NlV4Ur0aeWj40JWplJdS5aRTuPPl1V/lO4Aj0pBEXy4CyN4uVDUo+vch5WCh5L0UgcK1r
92lFzWqyLj3nXxYmxLNP5nLzowEj1WSqp/DAqNYCZpgrP3DwDLMy5ZEr1ciT6mqcvlzIFcRmrbrA
mBV+rF2bE6aGuTV7p+I21o73Ef+Qn9dJqZ6NmnDFPhzVxcbf6dko9n39jd+iFO4mU3F8vRgOWlTJ
OAbndP/Bri0H13QsjcmbcpX4RN5Wg5pifh7IE90iyqdPZRUt9xhJZcFipgeDG+3L8oU+ExGaincc
XfVOlQHeSUIpVjSC8qn2aJVqKLJB/CIuSenDJ2Y2y7EuT9vp4fdUmSMz44ma8m2B09uAqhYyToG5
+JQqFpxc4jaziYHUfNXOjlWnrCN2DqBtKYQ81bm5wPmZpQDHJxdvDbZTjeB1OdyUY6s40QsXtBJC
R1xbfFw0bKxs/JtyWxkjX7MakyMrJKMW0FkCcYh7Kj24sWX9kcDGBfqO0gQegNfApz/2QZ/lqj1u
ANYr/D9KV51X0/m0dgQd58h5Ovyb+s+hSw1rkEHrKoopmvbXtxfND1GWqVJWgpf/Ci/12XwjzQcF
DzS6YwNOwcwFtWK8Un/9l+pdpxFekiDyF48my9mKGHhJVq8J8NA3QT9r868ofqn2VLyF6l3MfdI3
3W8TMSa7fegLUcruqIgtNwkiWzBJRYiroDZrBZ7hEdoD7FSBMLEePdysWSLqaRAsk2NyQ2hQQo/W
tAeOMsMV3ANGymr334LQslf/eXLWBXevWAjmXTXNFkoVWo5AWR/NjnVZuSwPfIkLi/a6v10rzQ5u
VLf5oBNl0P7hBscpUn3erDx22LnQp1yEHWDcrjdm0Z64XV4Gg1EDi899oXT+DyvxvcDxV2ejFyKk
4OBhqmQRF2Eg8ltUN4FSXOw2I5TRzM3+x+3Q6REYSwJybaKsXAzRqvN9qVAvYbDlkBt5GHGdplY+
p0pa2mrW6uSlfE4a7Bv1AummzGkvHfDGeicvuen9dXBpPgmw4i4yd0M3vB0PrC2bgHRQC4vrYB3p
kIT+B/wjTTr8eApif2YfAR/81369QOVTPU28gXrnDr6ah1+pZFrgjqewei4wZc3MJiETxfVXUWHQ
XZBR62Ls12MA6+u06tgMIyUT7NMPo1fSogbgeCKZJ3KFHnW8q7HPOhMn8f0tPnrjfiMwlFOW1H1D
5ipZXD83hTxcQu1rhhSa9TuOJrso8uRi2y1wdsbuoBhyHYM6JkAefI4Bmso7zQ5PBKBuUW8b37/9
C+hc0t1oYPEwzis926laJ0F8sT1aOFMZ1pQg5lrhLg0SdEKaJFdfID/rNRsl+yWo0ba5WC594CdL
9uXcExZ/5mbsTf/bawPYs1Wyk8+huTFfYzypVWCeo/DPFrnyJwy4nCytLkPF42FR6eXQ78lkcXZX
GWwssM5jMAzd0dYHUgmNFg7AJxs+nVxNkN5p485qFRS1+thU4pK45nqHi07KLWwQOrswPum/cLRb
FaMh4EHw1Fy8poJ6B2kH5v3t4Bp/ysMvgCp10aNCDhF5KNqXQzQXUQ7z1JXmsjZbdFghkvEWNPvs
W3PzrmbYCJh8gcqWc5sEWJWqMPUSRaMYggy2iR6JHLaPL906ixajUydyMIgux1XAwB/OfO/QpdJJ
PJGJa2RXQQFDv4BMIJvccmfXezqvVOEDsekIfXtfZ6yjtSdyPz0EzfGTNK7sImhLGNcRbYNZsF2b
ZZ/6pUn72L2J6SeQDf7CpqlwPTOHL80AT5STkLJsWsuEGV21HlnELgMiuXCXit9IgeqRkpdob9ra
ZCP0Q8sNlXY4vNFwyZBv+M39bSyf33i8hezRwzUa9MtR0o0QKdS15XEE1NkmCVgO+TlT7SFLOngZ
tHS8Zp11hXYAmkZErouaAhn9g+BJQSci6WJpsKrNuw20Lq46UJgw+1OC7F0/AsWeb1NS8a+vlx8z
MYw1V8KKslKWBYD46NmrqxVFt03mgoR2cJ/R+ud06dTiWCNt9nIdGQCpfyqCOR3yYgrkkBPMz48v
/tOP7N4nt0i0za/hoayynLka4U+s/oh23dIOI2wAV056KxT7dHvJwsGnJNxN//Z2+c/B+jregqN9
PTLJBE1I5ZuSks5cocSf66NMygaVBxXxuy4XKqRRKyqi17qNadzbgcSoFpYsrdrXr8f2gFT7DX/F
XAZ+kk3vMKNS53/JLgfPMgcpeoV60LxcRz456qdOOlS+42BAlCRiNB9s3+W2BRhS2KH6YHF6G20B
9Xlwy2ovy1Blq8yPA1VLtYD3WoD1/y0btCk3Lz799BpGcuQl1YHRfAx+aoXAnIXThV8SRnWf7hwS
MrWZqkplQyUbkUtcikj2Aor/9FomG0sR9O80w8HuJg/8OARO8vC4pKCztLeQxOzvHgD5nNAQun2p
bocKcFEOHi6kb7Ov9sWFgLD/ld52djfU2Add4qpDCTUUbEUeaJ0C3wSzo+RgKLW1VKmpSuWhbUl1
OUpxE7RnX34SA0z2ogMgd1O+nu4mpTAC5sCtz1KEAQXMzYi4qRd9CFcO73vp+w/m6Rfbw2Agg2sH
/WgG1PwzSAb+dJuXdUh2xSOcWqQPx1jDeGPn6pMprPJYmxxHIlqocnO/ye76ckyKEjuDOaY0iuYK
lZns/1XI2r7C//DI2e5k3kTJFFiVv5ne17nIUYCaAXNNadA0DPiRQTu7byMk4HxTVuziNyzWyI9g
YwBflDbXtstCH+4lFXIjY68vFnOTCB24Ff0bw22VWJtMlZjcXhl7m3H5TlxzAvmF8Ksp5h/y3qE0
L0y5mo7cyCiz0TJlvlFexCDb5eqFlaAti/r/635R1dZKbucdz2AnDLzy7md6zor+TnTnVFEa3gc0
3qEg+5Kji+Xap7/XonGPFufdVIrDQMkWFaGARo4vjAK+DNumTkEUUPXI2+zhhqnAuz0p3HxyNcOt
InEkoWZuHEzR8+kSd+D8GduO1dvD5lRQY4qxHC5crKbRcySmOsaKgFqdyaH6+UkCkJvpFZOrVRQL
Xj54W3vDqndOiBfvQZJjtd9xzj+vPHIMcD0dj7J3qn+82SoQaWLNNWBdODiiQibvU9Z8XM7O6BIk
M5se4ddHhKcL6PtdWIjyIfJCGQbzMcXxhuC1p3LVbTmsD3P7OrvqhqJKHojANOFP95ZJ2lcCZye1
oFvA4QjepWO+gCTWVydf7QywLeV5HeaNULJsTjzKBiOm2LyiPFbi2q7taCqpdXq59GORzNp0qUs0
/aPLa4k0I7E/DfKXDUzXzSs4b9nrgon/b7k8SCeAZiPnHaHb7Nsk8MKGRQzOD8/JqXsgaDiqb7RK
ujkOcbxJYzdjdDr9Z2gFHUYHKsEbq6evHfd/2cmY7WO4lE4XIUGHVvZwE14/8YXBG5QV9k7pwtVp
MPrzVfkek/zvSiH8PwZDK7/Eh5tNzxBXmdKWi4pk93LH7ifPv5rM8ZB07Z3b3HFZfNZCcK3e96ha
lOoaWptkf21Aye7IQuykTxL+6+Pzrkrm50vkq552zZP1chToTWa1LEltgLz/GvaAHY6qYjXfSjRJ
QwreGXC57z5d53D6WNHneZv6I6J6Sdo95Y+s2Z5Jdks5U+J6lcbNGCA4BxkGend062l+/Kr3NT6e
pfpI4WDLpUkC6tT3emG38t9wDk1GU+rHPnKhChyojc750sbn24EtTEP6DFPxnN+DModUL0x5xlpS
FX85QZSan5UDo4vGGq6UftGAr1+5PXPD9akevTexjIEII2pw+8P6KgeNQ1FyactchgXWu2ay/AM9
IvzFLfLcMlxcbtlZYjD18w7mzbN1PZSOPdK485hUbKTkCtmDP/ORoTAP9o8wudrC7otjA5LwBYz4
MUEHINXSlGdYIhCpY0CG3K3IVnr8tA5S/h82udO6FIjXAzPWiU9LVKRCKZjbosKtcp0GXV4P8NMo
UFjQ9okHPR3lLcldTerwK8HbZWFMXn1hDqccrMc/xrJYxucz1gqnBILI6bJwgX1F9BcSXLYsk9Oh
rP2h8qNvo3BU8x7edRHSaFkimRqlcvr2fCjO2dUP1Pxf+61gmIhefc03RbgrA1mIDWhOxZdTuRTx
o15KsHIAX9oHDq5c0W/tVEB+j/0oUjvAal6r2cEaodDvhh+Z0xJX5ejueIRAjemlU9NcSobP/Ov0
3RmGKcWK2/lwmf43RnqoVrrFhrUcE15b+OuYAWKMGAHjqq4hpBABG+kv2crLKllOIODwF2alLfF8
owpLoeeOBzGC+eNMVIQerlRSoZZ4OxaopGqMl6g2emRv9owy5rHvA1N3B+6WaZXHuQ6Dp/eHbDV4
7EaNc77OHflbHngrlpJuY9zmxrhguL2xOS3SMR0TTfBf3x3nqR0wmpBkJfZRUNzRGhZ97QO1CWdP
xWofz0DhUYe3QFvOrf+KHNFsReGwAq0jKqu743pBeusaLvXrW3qO0/KfjlKuGbIQWMdbykd96pYT
dRE8/SdjoV4PbsEAWEPRxTowwTM4JaT+RfQA79//Msv2DRvaOP1U66z3qUW9lHOAHHecrLewe61g
bqrm1tDPSngl/IqeSMXDjDmgqVPx4GA7XDhyFHKgtxnSQtminWeN7KDl2d9WwCzoopfeOzSN16Kf
o25yHQgZFKwLJsgmuqYtE4YR9ZBLAEoeJNzWqLjdcw7BEm6NJaXj5pqBJCv6wfB06nV12op19O+n
GPC8ml7c8vcHbGyf8LsLK7mV4NXycbaGicFAKQInBbL4cUpkbxTWG6LR2SxTtQjq2V54QhIAmNJs
XtOZi/aCcCf2kV157yc8L0TMjxekwInVlr+fWkoNkuvAbxwl0n9y7OxXrXXup/6+Vwbd3TRfFbSd
YZLI4/5EY/cIy7uPkbGagSABmDvkw+Hr+UdWgAuUFcwfNtI+eDSCCtp0BSn98jSijUZ5vv6BJenT
lu4Cx7RAbabaRNPyskVb9XuL/tGr8VB7X0xEAQZ+8f9NYepW4I74ak3tb1ShmD5f/w/pTxdvZIHJ
nFxAhVTmxc/zwGoQX0UyoXUloAqzluRHBnUNPNL37A5tVR97+utBCt/oTNFfNoNt3+xrf5PH8y9y
1J5xDFCMg70isjhj5LbeRoOV4jGX6S91rxiLb4phCG4XTRbfrzr7SkKUC5+Kf0DuNdmroT9hxkiz
Apm0m7SdJWpwf8aaLiatl+R50dKMDPXm3JiUsAJydNR/hu4i8meVmDPcQ7Q5kcmUk6+kKz89d2EO
2vfjLGQCT24YmBRksraKKXyReUW/27p28QtsjIHO2br0gxK5LPwTnQZ6z2EFRG1gaw2wuuDFSTeN
3qmC9DSKKBsQ+3vKDfV7FBTkteW6PDMz7hrfKGW2yiOohMHhMQSo0HevSg46EJAxW+JOXx/zX/mI
Uao+9FOmzcTmDV7GI399F65UIRcoXF2v+7ENIQQYU8Nn34COTfylFgLKu6qe0KZOzAzXxcdIPUUn
lcOv45M/aBSGpiAM+rBY8remfxd78jLPPtqdXokyF60WciaGsIFmCQPvvYGrvCVTFCFxFqVFiuIu
qLznBbd4/tshv2RHd8lrOoo+sLEKXy3Mz7zwhSFbxRUK/qF4st9x+l6k82b3tTEVxrf+xVAHjdTJ
Qj8VWYCZ883zb+Jv9yMEhdBFSPBPgVO05yId3QULxiGDqvQ6OLkEcd3HCY6/+hjK9WGaIi4ZczK5
Ykcn7j0TOOTriw8x87rMotoPe97itWDBBdR6lgyOqJY94TNfivsNEUkw9vj80T2eis0ZVyFbTgfN
nA0Jq2AR24qPf5xzpkcMSwfwUpwmc1mIi5JsHb8j1g6tzpP7rehMPh0a/UGDIZiLWow7w6VwGCbB
VAmFU5f2lr15GYGsDUYOgHuLX0WG77q0VNwgBJmF9fSPLMT6tKtNw9SoDgSX82IOTQcXkLNYFiz7
/vbmNOu/o/7M1XysTAppz97iJzKN3xqp/+0h8Prf81CzW3tH7G7jdFQ3in2a3pSBBWtsptB6m5mI
DpqThQV0azvUylh/6jaEFZXQv0bXreKVMrV/8MpjVipVlPpNwv52PqzEkUmVhQuayNmJbPkJ7lIr
k07OOteBLQGfpfUKYPnaut2W2v+4TOaLE5qizetxgKtDDBs9Xgcm+gmtnmdpaS8bxr9N6iV2TigX
52QENG8HyEDu+jeC5vW/rR0WIQOZ8jb2tBBsrPUTSqWxo3dfEpBMiIvLs++iG1oYmHjLEIHrTXrj
vBd+zs3r2RuGBlHy7rf76UHaGYEpnNsbDrLK7JH4XyFT7A7lFuvYI1+cxkK0gGzoV1b20m0ibEM5
kKDr0Dk6nezaAcPjgeMa8XKi1JkCnDUZGKflPMuwgD5MJqG9lzVUoaRmG+wZGlmAGOqf+lthj4J4
I1TOEquSC9LfIz0EyZEynJbWNseEmAY6W+HQd5/2Df5xaClvCBPicZetPahZpScVT7OCmub0VWFk
nricUQOzW/pt4irM6J3WIx5QHWLJK2+PETdpaj7vIXcfjiYwWj9KWxkrmB3la/GvqhC3wtYKl7a2
JbP5xyT7N8CjI/41vldIRK34VHpwJr8DaQSsZ46BcrlV+EALCv41YrVSmYm+Z0zxoyWhLE/YCJ43
+mpGdnpwEcMI5zqlbXXgxxY382wjofiRBzteVw+KbFE1wijt4dAFh1aE9UL+f71Ero0zAUGGjFQ7
9zsgMlloIkuuc9dpG3h4ittYS4mTgq831xsqSOfShJc6efZNr/AFCxuTAazJS+23NVV1TpL+1OtP
MENg1jE/nkulW9ctApXXxHQdhaijF/RCQ/HgwzRecAUdX83sRrS6mk9KFPuI6+kEbk9kvffkwi2O
olOa7RhF8DA55Twm8IFHkKVjaHs+raH7lJwwoN2sLD+xMtZ6BPk4XiM/T3I7sqEudxRLqr96PNHR
WXUUPip/wW8qwPSJAFKGMOrRtVUCOn8VD3Je49y8t95COJmultMPBLGK71Qh+NYTi1eoZ8lOV6nM
lUXugnv0yDtHzIFL5Ff1/2vuu2nGc4LwvtUKRK9pQAWsRP4VhxGwVHrN7QUUaFbHJDc1G+H2DoTi
/yqPry57ww5dqZbYlpKtzaAKlLW9CtKRuYkq838mOiNKLCTLgjqvj1G0N6CCBzlBxtCTvMb0diOk
Ul0EjQjwiz/iS54kH9oUvbatC5tQMTQtY+T4dRkiwZdfEMqzLrYyAYdxpCx3btm/Qfi+by7jai5T
VvoTd7kiUr2TYcLiDbMs40bb3KIsAzEkQZYYJ/38F5oFphuhykIr6k40uQ65ZxCKFGxMukEtr3Yn
MDy/ybMyf/n9SIsLPgCo8B1EiVQhWGa1lEICu999d/a7sipMg1WZfDUP49FboXHPv2PbOBj5YcEl
THlbgooBgXtX0rExirYR0sc7Z6/6/+0sd1mJurXayul0StVMnTWKTmMABlifRvKIZW64fLX4tKkp
faLUx/NngHRT+XM7rZ2uO8hZaQY1faJ0lkj0qjwlMFLM6z5KNWGdfBKVBJqm4rZS3N9nhuBLa0b3
alWemO3PUuiLv2XZi0OVWY2kAFm6Zvqehegr6fDQ8nOxXpH25Lmq8xuQSOPFoOFDrdszoWhCYz6C
ulCkMh2qZZQMtrrFL18I16/PRw9R7omNLeZOk6W99RNhoQURGhaNADafuklJugc0rktMWtzoepMc
FdWXcr4hqmi42uBR7cXmDPUVtsI14GD0WyXpn7sCFxjyePh5F/gHIQvzL2CQCwZF3Jd1eXBLXkor
4TC+8B3gGl7my22M6ct5qiVDshaCmMKS7eiACZK9SVUb52yLBzIa5/eQ6uEWvtLk56CVw79gLNuE
x+wQVV3NOG/EMG9ofVeP7jpVelJ2RD8/58rUVizwpIel9rXSPBshB7EWy4Hpma+5s6Ze4eg6MR7l
cRUjAGYb3ZRCp/IftTYroqnntsbh0ud3vY4wjSJZ92fV0eZ0pDy7ZmevhIB49ZYH4kLwwVUXhU2r
y9AMpHMo1q//PpBJY1v98GnyW8W0A4lXnKSCMCTyBy99CWjyRts8RuEgHVI1FTSHgC1VtQo5TLNr
TWYoAbwaPxxdvNBaJ/tvwPEtF2bvhw3/rLWRy8rRDmDEcnMeBcc+jx9RGFjGfKPlOKXkVP/7Gg0B
xpM0JrzchYGZPJRXX05nMOwfDKojIjmIQabUMIJmPG5VlGtAJPWHS9CVJMBYDAOdkLRBBtSUr5yH
qZfD3tOe7xQA5G154t7wQ5mPpQl1TjsGfo3KBZ06dOhHdfjR17BwDnUfCwwStoUN7yE8uxKjc94A
9pPshz6Dw46FoMM2lVTd1DNGWqNcG3euSfe5z1ZOdW2LfeBgNJzCiUy/2zDQto+ULrAzNPD3X+tT
L8usumUp4LmlE3IS4DLPXjhvvxBAAych67BttLvrWMlcm+/sENRCcCk9dcBl3oisMvHgW1tYe/oE
DMM5bPHPf39L8IYLVo7qBHAzHwhL2SN0lH0sUHWmU3Ed8ANAY5ndXMkpJ+9bY4DE6/xPlY947yKR
pAZMZi63T3ouVfKgNA6vP1IIJhmr/VZVCPun9MZ7Ezswh6utg4I7uvOQlymOmlSk+29JywHMOB4Y
62+93WwZ5jwafTaylCtrWRRPY1AwBvk0YkhoU1B6xVelRAOg3EZ3hLjb2/a25OzrjrO6gjLjYSmf
XAHRdToHhteCUMtVKm/9Yj1U6KSukfFKycyMl2D1dpgvXymJH1fycr5/f2f4T2WzBe9NFZjLBxka
hUZO2wTM+5mQe3R2JwyBHy1IY/sQkSHnbU9kA5d5EDPAWRVBxDsyd+g779n/OAN2WXIWUtgQZqX3
9EOLu12dyrg0w1ArmIE53/paCxxUicnlfgM+k4rzLQIxbJ/JPL19iiU2BedfHRpHE93KY2eYQFnu
ocm2YCcC/cHwj1HC+8RkYwPpaCjxCrhs+wBS5R1457uxevQE5k6p2HEPX9Ed0WOE5pAA0PwVGxk6
WJuPBQdsTibEBDUgvJ6VbVMhyp6cgpZacftf6N/4RozvbNkY4+3m6vg3N5Eti3T5OiXv6moT5MOw
C0vpOXsjAr1F7JFTrOw6tV5/DrwPDnAVFu8s0zx9emzAbXCAqfW9icZDaKrKEAZpdCJRzHcJVE/V
ebrN0vLSu2TH+xojW0B8J53XWXOpCSnwRFOgF4VhzI7Tz8toLRkf0kD2AGAADS+7+u6ZcdvoNh20
sdDq6zOXwn2WP8UXqv+k9mq4Ref5uHH4vErNor/JOUIQNpcSkTD3c8l+S9+pTeEIpCF8FsdCeioc
iKTHu9QJaqC8aPe/ziSgvl05imKrjnWuGvGsH9SmlTtFfvxnd95Swx/qntdq2uuPoD5QCmA7VAdA
Vh/ZzH2z7MuD7LpE328G7qSM2stU22yCQ8hZ//sFykrHL5sKoeyNuQaOeEuI1xhWXdmtzpKqidoZ
0mjigbFU8MmQ5P2DTNftO/WznnwuBGLwc1Me8nLu3VFyGQt5qPsPbuTKwJJSHkTd0R/dmOq8VU61
Lu0y+Nrha+7q90TiCfs72+nI+6bX+EJYyMI4HIRXsXTVGt7QL4cn233RehHIu/WantnzD66ZMCLA
3eRTZtAWeh991ZWoFzJDN5gvYrIONrsbrsmV81OnxfhtSj/ukr7gjdKulFRYTxTaGIKP+3jgPUPX
kxeNJd5/lWzFXzWp5QBYdGDVWrD9C1oFHk4G/4CdeuGFhPD8sUkCZ6G7N6F4+veyqyfwBWwJnsB1
EfZU3iErq/tmieQx5s1qlIxeXvoYW3QMh8dEWGrCZZFMsb14WftZ5XL6nlbVIz9X5Pzv4iKyrSjY
AsHKI2ytzzsXXH7kpWyEsK0pjq6q+ZjQTL3eZP5dygNo9n1zyZbrdaJ0knKk5lYivSAyfU90cTKU
snhr63S2qrSMKGM/GDGd/hsSo3RCf0NfQ81rnFEwcw5smXwcSSh15DbxXYhl7Dp8sOcrIWtNoBLJ
snJd0rBJMKQY7eMmcPnqpx4DQKp8GYYkLbMV5Vnca8MuO48YTVLWE7nWtHbwir2OFr72d2XiJwAB
c0UVL3tPwBOaYHTXxqfM0e+IadU8d4pe25tQuAzcC+oeHGRXu9Ce99Ec583cvvZYZWoVujYGJQPl
j92Xu5KCex+pNMHZEexXEtXaKa/cxPU4Jd7YdhK017CuHg3MBiOFRpDmFi9o8DLgyHSXGhuha5s9
amkhtH/bDIMsf0M2+3qs3BslIWsPh4h4q+H/o0mgyYXWc6jA6R6ODfkfgomExUZM0If6lrZoSzNu
mBNzPt34taVo4NBgySYnTzX9GJZaEFsTjlfsmB2rdq0wO+ifhzE9XDGJA0c3WhwlVh6PVoNIi5+W
V0wIQ6H4wYk1yETL9STRwKD7CJzeNcnpb6R5P9sGJjcxYAya3oAxS1oMRtOTCG4f+Zrx/lXy37av
5PzYGt7uPlQaSum2CSWedwBATR2flFdgV+CCEVBuaxOlXRmxKiscVRNnq4JRKq5dqlFpUsBgN/H7
g5esTfZNVVkb9o4w9Z1tvAw/36qVo3EOL9gS50NYFzR1yV/0u55bRMKcG6vgMQ9IqedXqLMKQmyx
Fyvw4nNV00J9n4gdV7HD1MKCkWJ0FSodQrVmB06Hyf/5GV0ECy7cKyq4zvtGHsMPclO102SQHNYj
cc4bwHobToSU1qomtYLUdqO+RTSq6N2SEWyRegt3yEVMG6PUmuwGsMmi9Iifvs/rQ5fStpyUxNWC
uy0T+PaB4Nf58Y06WQJxgxh9PPpUTDf6AJ7eEkn6MEloBItMQDicYCZb7C/Yq3abnlv8VuITKlDw
u3Z6Dt8ZenSfa/dElPa0ysVjToX04lt4Z47aWeIGHb2EFasN3P7utqXQDputTOUnxN2WAsMCAcbK
sSIu7J3DnqxzP0KamXIy9gBicCQWzW3fNTdgsSXFNmhfSZHY2iElb/gPsJZG3QZDGNKaDXyoIFuk
GEwhvQ+XdueUeh9N4taCDFSyb2FiXJlqI0D3/8DWU+IY7MLJCY367gS4TKrUhl+Ck2s+W7shXBQL
i7Zehveh1hE68xwAzarfMpFlaYBeuiDo4gWmNKSABddy+C4iT1eLg7EnNPqvrghz/noZJwHDOKN7
voRj6Am/JNFT+13bmp1qw6xMtyHG3r70JbS9SrUo/97/JYhp7N3UspDVUX1uUBs2jKUEUfIEFXaa
gPpKn7LtlYK4AMBD6b0GesHMo+sdtcRj7vRFBKn4HGp/20lrz8qGhORVIQuDoe+sYe0vMosehsFm
4s8A/S8voflqltndzCRY6JO5ZlGBwr12Vfpq0Ub3+aMVWb576KDPFCsaSeizJ3UdXDIk48a/NEGu
Ze+UOo5E/+JJqVzFVtM/ypg0W7FwGbXQ3A0UcFeDDR70lNFxgd/l5u+kTCD6Gba7jO8b4jArqYWj
wXWRrHqkA69BKEoxPDHcdGiRN6qlkfbN1dq12zaE907vOJOTdjHIoedP3AiEyHEjo7yrT8gSdYC+
guGu61uCFx5Veb8ft8b8XUxYHlfyvXIaIMIi2zN/xm+yL2SFnSC7E6qIbOxAMS0Ua7gLrzLkNVHT
FwbF+9k5ClDJQL78FF4ut/sDsNFmpuJB7BEYw6LAalGQtzEs3g0T2qv2hGosQowBLNHGz6OshrcQ
o/8aB0XYHgxYT2s1aeYC7q1nJI7sHYjqDl34FVn/x1LjVlE4sqeeB86K1kGKt8Pycw1/R39+I326
goQ7cG2XA8Vrb5tnVG3OtYcTwno0D+mQqpm0GRyiBmi4JohgjR3+4fh1+qght75XSNO9dIexzvnc
ZaA+rFdNGY5Mnj2aE8q1ceUv3UdOq8o6AlXUTWFdBw5iRhX89OATPanzuqwJEuQCCS6/6cdWsABM
EoWBKUF3BzsRR7xEr1yApT10sg1X50EKB8quF3LTVShzFu+8H2W7pJ3IQrAGrRdz9BoAyG1QmtlU
NCgl2aR4flFaPYpd/s4mrJ/VaaGgYvcIHcKMNV8gMNRhf9zaaTQTDALWjPbYo9IE0CSItnKVX1M6
eagkiFSSVeVi5NPQcs+ZikgXMPxzwnXGXAJBBY07BmnMN4S6bMM4jOtYe8igjNzj0Lg0E8vzxhAU
IjtF4GmNcpwfZyMzX7dGdtmuf55Dd4y8Gsv3DwhDp785LobIA65A3YSi4CbgORRrMwAPF7JgIr5I
SvpLZbxDPLLSfTJxGIxXDJt5iZ3Y2h2cIq+iGI5Szz7h65cvtGQmhAmxyZ3Tbo3z8iJBlO6eni+F
z+pqKjSOqoqHnnAyPO81rMJxSm6i9JUSfr0K2ZDfyP/jVb+zeFfXrq7H7/3HI93b1BUXxNPoCmX4
r0OWH8Xln+fhwMAqMUsFJPd1aGLKBuYuamFihVF90HjlewltycDl6fPYTnLwZKygiiuJ5yl7bKD5
zj76y8qfS8GwL3OSwrOhtyLMmB/+yqZI4MKponU+M32Mnspug1LyLwshL0A9eYfrqWMGsvHx5o9W
OBFRhtuDLma7mkbb65xBgcPDDftYb6afYkOk2apukINtqX6AtjQ/C4rHbUdX/tqc8VSJLy0iXlzT
MqAeuFRxLHWrmYGK/wynA6rEYJpr9N0EXgS5jYrF0Vp96BQfQEzoei2+ph6cg3mbMmj0ma8HvIlC
yX/HPIQO0tRIyytqYAzYBrq2HtC9nlHqhq9ymI1G0+RnSgCas5y7gmGm3nztUC3tD07o6bF3mACQ
qRsp5r1DYxO8qonDQIdS1sQi6moqdfQuYmpKT6ImneyYslWUf8G+ZyUOmldP7Mn4KWaHlNfabqTk
GGwWYmpISrIonpuJfWA3yPw5/iEKGYw+U/M8qQuGfKGAKegDBXHD1rnuZNSwoey5wGgCkFU/3zrJ
FCyb/uhrMeQLDQ+u9EdSTAL5HKcfBJs62E9g4tnnaJquC7zQXO9duUpU9t2KGToRFldF3TpIB4LW
0LZMSw5yBcI9WBY7PLrs3iSY2ppqB2GofrzvM1U/Kgf12Z12lf+iPXJB12HDdQlPRcjYIsnHk8w5
oQ8LwoMrFTojAtYeWu4QBqh9RYmh663q7K+mMTpcOOyHaFL+/zVJ8+83iuTrD95nqmC7VCZswvAC
tna4bglj/kkWCau9mW5vV+qn589PPpHeJePSlQg/ro/E49rfKpjizenolEBVoXXhSaTNjIlrGA1g
S+VbB/faxXPd7amSLNvEuSveX84i8ThIXSG9cQbuaAPymJJ2ympFYM80RHBbSPyMhgrr6K71MVYX
ndd4h/0h92PMzqNNRiotDmF2zgcf6gHCsj1wOgPXIbnk/dpKZvx+b/AKcm7/IY7N7+gbGgUyAWO3
O6I3Em699nnoIO6tvphS/KlsCQLmLEX92fSqvvJwG9muMCooh8eXXpZ/5JnvRQngDqC/lP9FTcXQ
gC/DDfzyPtjkkPwAg+GypsiUON2nJJHU8ri/NNP/okJ5VGG9+WPGxpnh5y0EZENaF20YdqK/6t9s
LtK5AH0TQaDl6jv+pbXP4NwOeC3xjBCLCpcU2P35sMRIkvqh42CcDDuRYm2M3WI8tDitYLNvTTgg
g0we4oweztOd3kWpzNIaYKxZW8o0nfPFThzUSULIUJk5vBq6oWUeGoEL5Wh64zHyMLts2qvBoPNY
NPRkEIfHwKeMxvU7o3H37aHDls1gNoxbar/47mURA9QZXVmbQzXhBF94OT4J/46TN3olFReo0owG
Cy1cqPvqnYR3sb716CuNtZTpLdLA/aBtsJ9XUE4yYad/0fDHH2dacYHFHpEOStJB7NRRQyHpZZZd
UQfJlnf1IxNmPa2/cCv4rNSGyfOh3ScTo6TVSOhZQjL6+BzayXbtjMnBcLM4pEOzWO6y4zM1iYwC
ZXCq7afAg7YRmW+9/RhGdVtcpXFiA2VMylP3wcRTKBTha7kSIBhFUcvNLhyWLXkrsjpF9997F3yQ
3sfA++gyn9oocRBBXibLwDIYhyPh8q6q1o+fUDbrXkvBmSNGAuBjyOahsQnlS/8kmodWYNv9DCLI
oVnQpmHK+zwI99PJCi1C2lM1oBB3z4GPdfAZQgLWxvS3/h1G8dWYbzR/rwqO/Sv2zia8vrao3cvG
j+i/4nZA44ezbzBgqtoFz07M7utQzb6IdauZCPxgPRuVDIlUD+EqkUCL9SRGjrf21GTbLnT2k97b
tCxiAKGbZ7VNfFqxH8ES7Tu/IcqliRBJwy8bDLMHRX5YDsURPDDBjuigbWmJpIiJ+etAwjveb89U
3R7V8XweT4l+MoN5TKfz7+n/JsV5vohi7KX9WqC+fW4fZKlnxOaep4EUtqrmYDICsgJgUiRxWcvo
Xd6N7QZ1q4Df2NV/lrRLkEhOi4tQXeTJtY4AvQwcbIyR7OeXBDXFa/06mK3jXRM1MOnaQDjn2PYi
vmiIjZuI4+B/TJCynlNEqTni0OyObICrcL0ATKMIaw300YT2VamIjKbNx4QFXBwVRcu+7J9/e6U0
Ao/u5vvVLRM/G/ucUTSfMO1vrspYmwApWXx/n6b5HQIXugOjPUAGyA2eALO0pp/j85Rk4whaDitm
w2oYh3qbAfigBLVJXDPySHHlJvyE0xWVzFMs+oLWDw5E6cWyK/URGj1MnvealANGSfEcxaVg/neU
sXT3veUmD0n7lIySuNsD8ahEhQTYLfEX5LdshcbTZBQheCh5KHepagMp3k3tWEqZyEngfzIQqlyS
zuF2SdiwnekalsT6m4HwRXCG85ysJ3pvjRND34SlzH2qZjTTmtXOpWq5ar3L8/cU3yqs+TQazXDn
O80sI6M2SIeoMgqX+W+SGMKHDs6pJKKcjlkqeyesLnLjVq0tg+ESh2c2y2H7rN997N89J0S2aEUu
HPxMiCF40SoIxrMlihrdE2jlSj0FTuwSv8TqWzK77qbDmRctbJCuaWXkebNE2Q/8h8QG2p7Fo6wh
CatRkW9nvY6KuW+OqzvhLRVvLWA69Nv3tF/MuyI7c4fnJY8V9ApzZzTf0MY+jdl7AoYYif8FWtkg
U9pclETPFW+otfPblrrqxPWZWOqjBc+oXIkDbr64WTOpxY2c2g7h6kPmaqMI19E4UXyEKsay5WGY
LnQG/11D4/v354bNTbV5eFLonD+qC+x7slM28W+4obSxAFOhplE2dnh9LQsx/xefk0EijYIk7oxE
re3lzDQGn8b+6bcUQNih0UQVLgAYw2mkvZyg7GXDxucX8un1hij1z4Ew7/cWEM4xgKS/3jrQQNTE
6XRRnDXOcWy6rTnQNXb4Hx2nRqbhWB9hIo+8GAPhlj++G4XAxaKvdHHWFwlI+Btbd4b8urMIh0h/
yFaFgDf18RBf/JfcTeho3Xzs1byDDJOT6r17DLsBIUfilUtXH+Xv9p9UxYNJx0f7oENFMbdlWudL
y/kqpbeYkOLx593ZEvfZKVGUGvzuNAjjoaU3j0w4lmii5RVmrjh94RBnZLSPtM5rLnOQGXtPTOBz
/KUs9D0GjhHRXba95flMUEuZC7PTvnLiQaqzmyqCA9lKI2FJF2rMbbONNhi+Ie4fKdyqKw5EWhE6
0EVgWFpQ0vtLD+Y5XHIYMV1XdRpnRlv5tBeE9+WZJjiOYsbQc5JNNSApEozAfG+etZYTcQJ5YVAd
MvivI3MdOuu7mcWBKWlRlProGkGwv3dsWOWVro6O8ASb7zbt0RDeK6vOFNwUl+/XfIh9HpIeKs3c
YlqmCfGg8RUi6FP7iTV/ly1YZxMS5JXNANFeYpuIq5hFsGVdpdKrEh1KWYB7DUPO7Rpi1u6hFTDP
6ZN4OfFJ1wZUyT3Fhcb8qj4Er4lpW7mKCrEe18fKwqaXSeoj2Cavfa4dLu/qCWW24Hw74TM4uqFl
JVA35VuMxcmZWH33GEMrGUB03w6GfPVy8276pHeyud1D4LMBkZ7QNE/OcwlNXAWrhOe1BVc5Wzpg
XhDyX6o65vw5qoUVV388+3cJicHY8q7MZXkkLTK1jzwcfGGbVYALxuq/Y22VxYEdz1SSdFGaFzdq
/fG76hn3PG/IsAa+5H0gTe7HorNhfEngYvYiM95sq8f741ET9rADYAhn7tzWsPSJ31drsd65qGJ9
7rLwSc6XkQ6taf7OF3bXVtQlBGSIDrlJiDF52wMI6ZHEag4KQn2FYkGYxqZw9JP5sUduWoRSEFch
DproMsGyw1XXOUu9nb1USybJTAGkiI4YGBmVuQdUT1iPkvpNKQqNDR2/TGPzfo09utpo8T56m/Cm
iHZ8DJ2H95qiG7TNzuosuYcqPCLmFNy3R+Qz2REkSeb+nVeNu04/FmL7T6JYKQGZHxQBPJEUOLZU
3GgCSOEsPHbk1jR/fzJWxfDpC9UFLTr5rbZyp7g/18ADtXSSBEK8jqA2AZlYtoe29f7gHPr662KG
XhxKkcaQA6CjGrl5vpdht9sW5w+7dszI883t8I+X15LDlYX4CQtKQV0tbhJaE5STMEB1RFydp1lf
qh3U2V0F0sau21uKyxIGQpm2BXAv0nhlVKSNb2ErPBRrWY5Ko+6r+M/hAMU2oRcfU13UWm+7FrB4
l6b1jazH6dFs8wv6njVLTEb39SE+f0caU7qa/1vLFW8VANbBI8V7nWnsV6zHmsWF6tfykJBgRqve
pKmojTpauzBC2amUX1bb8GtxHvzn0rrpi9jbd2vv5UK1an/dH/Xe6jgWvrBKSFzQlK2C5UdbFYwc
QT8rztTAv16lz8bIZiONP5lulDN7jYiE6duzgN823f+wLragm0i28n0BDp+KZ8NqgIKGqWiegE6Q
G2V0mVSMFntBiPz5NX/r5NEtzmePhSVDYns/w4MQCbs5jZmcMVRgxjZoZL1WS15ITfl7J9ps86fV
h/d+DTABYVFtJwQ/4UJJGw53WUL12TFwNAijsjnvgZN/nBprGZcHg1nlCnmCC3EC3P+U2oHVei2g
8mkR8uzvzWgd+am+IwAVlB8o7oXDhsaRfu26qtGItQZWtOlHCEkfRGheLD3uVsbO60DzH3vAxB7f
l2NpXGLwaLc8Y1FbMX0Tv9BaHdMMsvhCI1jGwoobOUjoruttirARCxsiNyW8m/hr4dYPqHEatWpM
LUP16mrGIPgQ7MyI5jRSOY6gzAdvys9NLCagbPtE03wcdHCAlSccQdSmXZ0CV1R6ZiaRjeMq6xys
60GtG+PdDhQNEbFOM4dkp/7ispXmaHYP/ZEnLVCUNz8xVI5L4NTywxD0drgFAuN21hhG3aOzJQNI
EQnVk4oawhtfXMBOMWV16Oleu9jCyvIG7PB4cgEw+vHVVKTYiJUGcf5UHVbGKVe0+MhNeyIpEBZO
rSJjqCrPgMt7m6SWrh8Hjglo8jFhgpqXaG8JUxCKTfvtpn33e1xCZpwx6yBosr5cLLMZJ32D2DcQ
4aWnWP1o6kILP6g6rabUdZJ5mNt9FU2Y34CNq5iahZg0CCogkLhJEbzEnAqGdvjvhh41JXM9jIW+
iYZ6pzoszRWXQnZZ5lHDKHLr0i+3pE74WE+G3R4kDEDIUka7QEIHD3MyHnjpyg24UQp06sTUrB2C
Qfx1kvqYi6FlKiJEIBPA30Q86UYlKD2Qiywg37K5pp/Ry+ejSLn6gnrYytjGGIWe/5N97KWmJ0wP
BLFo333GAA3Yj5qCdLms2npPr07FhcyzDUWP96XQJs2M9Tcs5SKrkpGE/JtaiA1L62/8eGrLRsi8
fIR2wbWBNVxXKrVlNvPV8gGk91kG6ewOL4heKw4X+XT/ITypC8v6OpnVAsE4lKpTdi5CEEDFkWxn
szIApP1onudvFkbRd6OiNXYcRfdwfY/K//pVnAiaCCFLpobHAN9AUDwv9+dceLgVXLb7ZCPOhNBy
3VcjKJA5KTTCGv4kAMv662usrQ5xB3SVyrU/jgZFhF978DFbcFY32SPYgnPZtVE6b1pS+VJqP+0U
o8NvQMlKCm7L06BpKvxB76uhQdHWLPRI610E8488YUsLvE7cs6AINN1Z8bHPURxJZysNW/wIUl88
WxtIEKWPhEWWoOhaSJkFT7GSQbMCNfirgzMjxXF8t6msTz1iGvEFExv4JVTXVcgmuCnxUn5zLY0P
ixfrKg+gaDbtGgmC660pThqFLTycYtux09iq6qsO1bbgGFrMH1YnnySDAjQkExsBKXLFCcQqKzjT
7zM9XSYQPh15JF9594wsCt/F5x3qr9W69wQe0+k4d++uyfpkOOiHlId5DYCU4UcgfkehnIkqcxQ2
uWyBhTeXSm/d/3KKZ7DvX6Mu2ZDPTr4h48ZFlDbNV3WwI2pxwXxwf4OZYDtr1ZckiWF5mK4AQ4/a
rVvtJAT8W2pIiOkhWghHkVa98wCpBqirs2YuEWWWWI3zawQb2cMl0wzXh8+Yy+Ri7bnRfx6ex9cB
jfV2IoGrsbsXKpLWVd6BIq/ENj58qW9v//d9TEj4EzThkC8zwZQlehMeIQWtjA8C+5b/jph4BqeD
m2qtCB+MnBdhqXc6kSPu8p08E9iKhc8aQBJxNk0WbPBBc8CXQGyJAAH77+llzQNWTZkIyvsiTUB1
vnLUxrgudWWch1iiTGMUeC0mjTi+7tvYiUMP18XevENph090rfccs5a0ac83ti0ex/e5+l+nF+Ew
iuGW8vjR68rOIln32QpE/BPN3XUF9TxiH2xf4/P27xlAWRdx3+Fak9DC8b6bQb53SdZmVA+mAQwr
Yf/kvN7ER6+OYWLXKzLJhtNXOvG0El5FJNhJyAHnBaAG4grAfavOmgBbkhtyHn7E3g/Kp+RzFIMO
cdn25ew1khgabWuN9gS9oAJ+DSxqfZJX1dICli9JMwQf4iBH2m2Nlt+60NsMFqsILgmGDDCA75nm
DXUadrjSYflHA8j2eGBYXtebmXs8VINeVi/9PgklDt3ZKv810kj0Izw17Lij8lWeIk+o3hzfh4n4
2qmcFB5RLVh39g6OBYShoShaLBQQhBrEJ60Ugqo/FbRjBgtNi0kkR/eh5Prw4emboQzAgmKOO2VY
RJL7mReZkQ+6FvbuyxkMeHyOByzHletvOdjYprzptkJdthT8OyLMLBBo3sfzoHV95C91PGP1+kBD
edG3tXnzzMlgrZMSdOjJty6Os8C2IN1lQxrT0mdXjMHa/RIxgwUbz6agimU3OL5OikNsnjkB9CdC
fSe7TxSR6GpEPCIjhfhFkMNeL5M0yzt98ZL5xwP/IsOLVQX6EXGPvcCFZozzWXeRC1DXhzQAMjPq
L2+S75zxh2/Nbac6PqGafM17N2Az3v5OEkm5A7nvtOl7NvMgyeAXzzzUcLrmSbxhai+pv2nu7qVY
2hKW0/IcujfAVxITURgnNvt50I+2RH4CExG6pQxN8LlnPHF5+TOf7Zru4o9UOuer2iMquvr9edR1
Hhz2J7viQAmt/ufRCkzT/wUFoNGixltnhoI1OMiMAnjWrL0XCrcAZUC+hqK/ZXrY8G6MKcwZVqxM
yIPMjCVFNJ0atKlYYlmcr6dTBMzJMs7uI3cSf6CTdnhHdZK4ICgCuWIB1SrAcd56eDNWxgF+430H
4L3yjn/o8T2D9QpOlZ5+6CoANfrcFO0L8kFJkjLamY/8ZoRdzZ2IMiMzcJ1WxQsxJeGOnupnohER
rtZaR+XYKVGON+/AEopZd1FuYptRmPxVdbQnhCw8i2aozhQJf7zIsvJytrXtzQjHzF/mSIHXyYhC
0Vk9cG2xGUoLBXTU51+bd20/cgwGCzaelC6q/z4xeQ2ucc4KxkNVCPWZMQqqaf6EiquiEGpT2nxf
UkcVDJJnAbtehJixHNDAUK24zdXZMP613KR09IdyL9xPNausz3Uv5p9t3+kV6Zfsexhbrc2J3QYH
D1BYti0GYB24ckvKO5SfuJTX+/iGGzndqlneT/VcRITyde+KcSB1EojBv7xdddS5WVD3i+5+xTAK
6n25CplwgsELaPlCtBz0JbDHnYMTu9r4WkEbFsO+Hhc1VOzlI/6bfaOP9PRG3GZpyP3Mns88BLBQ
j4y9SRWQUr6GHFIZG3agA9NkCVnd01r8ajOq171d1y3J39iAcO5jCauJCBz/pxP0vI+MdLG4uot3
98Baj/u8fAsHsGePrTPyOVsmL8WhpI55apcGrdBEMKDgQKv6By52M3VoOaWs2fA12PYLit+w4tJO
2RuGWH7RiRtyHIJOCYfLmxzIwCm0EzQjbmcT7D7z4Gjzwj4H22VJv2ihdonfA41dVNfBTpRxVeds
Z1FHWbp5XYUNWC4/l0orkbHZndcaHD+wc0XnGPrjXYVINJ8ueYYsy3XshGV+C1ObEMJT8Pxli0uS
DBeZZQgy5tGO+RtMzc7PebBFLOnujAnHVzbdjczX6JEhSA6B3atYqxedYIAkMn3jPg3rUJalw4nh
j7TJ4uNDBdperx98zk8lNu1iwMpNYfx34DZ2wDALrXd4Omis/G1Jn2UoIiBMYMuKYVHciOymSt6u
vOKiqy0JW6vxzKt7AMDsBdw0LfoDB2mjldrLCcvRhk2wRG7+lMgQ57F6y9GnpQxcgDTf6HpSyGxq
ywFw85JNNO4BQGd9of0CX+XW3re3tRpNhMexCld9DJa/nGu5Erp62lWqVm4HmZwqU1e7W2ZQ1JU/
DAuUIFVkLqUjsHxPb130p9A9Ywc2XTXOOphNTysLHUdwE98YLZVXrAMTRrk3QZZBb6lmPxH6J3w9
6k/DUAdZIc99WbVelBqTSusPFXdNGpkkbmax20TB3QMA+weaROUFrrInkwvBJS7k5kb8zbQedjX+
EcQD7afp7U08Pvg0Vsw2IfRelfBe4lsgZASu4B01wfjZZBQXNona+x+8VruXt7nmxGQr+jfXZMXJ
OAksNBxY+TCKKaEnNTzstKNLab6y+9AQnbKIb1IudSN40tsdH7d/uYBgpnsF+GT/yqG58z/FTuaF
CkOqTrcWZ2JkJH4PGyaHVNGb0XrPMAYUHfrAJS4blmS5m8g7bKoYb5B00xzm2HHCsqQ8S7/+c3WH
jS84j1un07UHMwLvNqIdiWUYVlr97JBEY4CuMSWCOfoysejbEzjAAom4vg73W0HdEi9XOEU83MAT
H1RXhkNakaewjjJVLrG508Jy72dJLd9U8jDh95pTNAChYu56Bvya+5zAYY31wxXUPEG8QTfXym9O
ToRGEHbOiolutsuzHoipI/9PPuE3C6TBcPmZ6dnRupQ1LGEWhgSar4F/tJvhc09nhaVlSW9p4K5r
tgx3uvrEcns2BBVLKzQSlI6+8EtQm8o+LNlJtvj0nDrilh+8nC+kbH9niiL76y5Ks9od9pM3I8Ox
w16K7DojFdjvHGT5Q23dP57iVfXMXBsBKk1rFaL/FwpWjlIyMU8v8B9AQEoj107/YS7wAh34SSjU
+ezj0f8yrT3BvOZSrqWD3eJp9bYgxfpRspZf70HydhB+VpZ4XwMM4dGoxSgEOu0Da1fHGa1o8MS9
JblKXvk6tx1ZPS+H+WQofKp43UhbJsBEz6ea1O7y2EevxvN6yM1pVqUaPhmQtsvy9Gq6c984rjRP
Txc4oXetQN4JmHxqCgo19DtFrZBBFt9u9w/JIJ0mdT7QeLM+esdGHljMFxy9z0SxpGsROYzJrTT1
t/m188aDD/jtrB8z99seLlkAtZ/9DjWXjLcyLd6GXYIP8rq5fCVOB2WcpdglzL8pNuhzuAFu8ESK
FlqWVXNegZFn4W7MqCbNQftn/EMpxqFGkvFLFgu5p5uAY19dW4rbIoKjU88jQsp9WNIJ9ECBEleS
3gOMCDa08lfs1H7Vf1unO9x/aMhXv/skXOF3Lb4YJI/4jIOzbbDDS2/uj1rbrKxRG40nrUjtbRIq
uWnet20vuYuMq346Q+cqizscwLJ8nKdcSO5ZLvfpUidibvSixy9sriIwd+RK44KZ37vznb9x35dA
n5eazMa85Vtc/lUHDkmqg2Pne61oU1a/EHTZieyfr+maApDIVk+Q3FAIH/hpwtc/pAWmwh2CzbJw
l5hidVGwVRemLEtim3eFmNU70wTyywqhi8k/izef75zaxeVfF1Y2loSEhCQL+gt5IVm0lunaRRZX
ntivp/2GDZQFnO8BDDlpSEn9Lr4sRXiA5U/edE0d0YVQXAwsOXU9ZGbQEWNYsMYKcYdQH7vBTsm6
tUlKWzTtVfdkClh0OttRJyp2nwro4do6WcLxehxVs26h6JtCNmjcB7vOcYK+9CRUF02pbs3uDCXZ
uIFvHsec7eHOSC3HJ8HHia6tIWBGMp1D+nCEfRT7ZzgAJa+PkHzwKGli6PLfv4JJl3KciPqOr+e6
FzQJSBJ+tCFsT/x0+htd9RYNXPw9XxddA2e9LVPnnN6T6UitJ7YWfQFSvLyi7vTp8R3sQEDcYGLZ
Cz8nKKZWxxzIZQgXCBrCoaz/lOm0Onp7Lw/fb0+DZVUw9yJsx2pBMJWtVsuCe561MNljYv98bGWw
HdX66zmQ8430qXGvX66URLVCYlXvBqeEDEn2ZXaSZfXnIwnim6C3D+xJc7Vrr1h/c577E7/yq84U
UHU7V6wsraYsUTDFnE98u4MnEpn8TJXVsCWKTaLIjlJgr3p+jDckZ+mWQp8UrJd5C+L7zMEZLGG0
/tDIzlO32IU/J9JFw0vGpZB3ZOw+hB9axo9rFlh1nP6OyFYz873BV4kcKRuMs9RiU4hbuPOqgUmO
MSHfAD3GutVnfY1AjZSuV8ElyHYjQ7GkAmCOz1kgi1o1bb0lIEMMiBsnJ6QCzXBzzX015ZgPaDuD
RLGZwUKNqjklmgClxxqo44dYKZd3yGnVQniGFdMj5Ges83LLV17nZmMV2VkqJoInT3xx3JQflwZX
Zp56bB1C1fp+COuhEnVC5NbrDxUcjzXwWrEkDbPDkAI1gQjZPDZeZhbGlH1Qw5WbmhfFWaLChnhH
GMhEY4n6TIIsflAbFgiXJnc7LIFAZmTXDnKb5bQZoNVaXShyrpUJmq0VKLne/Rs2z+UN8GUOENLB
RgEK4ewkLKoLuf0R9KrrYOyDUVGgxB/tFKWmYVjN6fYKQ2ocEtJU34d5VWdOx9S1nJ7Aom+wEC4D
4bzxi1/Xnqonm8fR0J84sYPs5+16saLyq2W1YLJGCFmY4yhmd3BcGgP0fozuGFY8z37L1mRKP+j2
sHVQ7jMG6/8v+0B+dRm+e/3u1NpwBimdhq5j+B/a7iMf19aVfjH2tut2AKJjTS3rKvlVCO1cMjQ8
OCnypiaFgbl+cMxeMri5clmBt/8yJ2UAQXfCYXmiuPfCgJcz21yA3Zj07PrqL3wLKNQAyCsa3v+Y
MZGoEdZT0MrXplYSemrT3n7c9GrzMCOyewrfinfGZe1Xh/T/oJXDFAiM7rEvKYWDQQF1FDJ82D6n
hdGn3/Qg/PB1SCHqsAkXdfBTd2QXPzhYZyLKNzjrks9dwkaG4eqwkjtve3QVtFiL2FjPV+cv3Ia+
75xE1qDtMixzXvRO8qbviyw+mwoopxtbRyt2VfKX0n4d3tC2DMBkFdZ5a9j6kEPFIF2o/PY7MOiO
FEEhWfTz8MmIvqfRaPGAWDmIlG0n58G9F/w0A96fjPLJWvN2rOJG815gwzf/a40TwJHDswpw1+HJ
QyL/VfRUGb98Wxp1q+WAioIm5ZXWBtq2YAoVJGTCRlDl2mWe0pzJanapjvFLEXFjTemwa8YRCev6
cfK+T5yDuQTn+ev3u8B5d7yzfEe2hmupTQZjv8mZ7HpkyHObYdNOP2UnE7U4+I7XzOg3CKgN+MFl
BpmoCTpdTZVh+c3yt3ctoMDtUCIG4Y0kzShGYKgkfewjVBhABDpTjcNj4vG5eRY6ER4WowgQJSIE
Ch+vc3+w/NtXd1F8Efvl8qfesXtLXoZRvf0wVBZU9oB3U91IDXNDqdfRRovhUpigCj6FREkZk8h+
6f5wpJioxTpKPgHYInGNafjGTVSWZ2Ie1n2Hy0Q6zMVjUrP/dGUSajzS5Ot+iAZVP3IlNtjOUaUq
vBAlrdiA9GG7zmlhnJlezKAJqO8Dce0mH3PSZ3T9O6SEF28cK9wdtVUR1iBqQ1a3MBJCV0abhVDa
WFMbgqIQljT86c19ZDaL6+R1NZCh9b2B0A0QKmOOoeNbctrpuwkI6juyszesWUnOibYCj0jtQr7J
+FxF3T2z4uo2PJulIV4hfxSxTpaJdZKRKf0bEwkeAFnfJtbierdGIxSKb0WjX/clDvI82WKSgMwx
stakzjMio3fqLAvqK8oUFl3j0NeQY51Ji7Czr9BAmhOCbLOtUR2F0FZAU26TxAkwKWVMtA1RB3yQ
PkmccUhbs7x+Zdt9oGBUW+jvlkJ00+vt/tSNCo8Qa05p3VPoTkeCPJN81UGn7nUO4C1pZF9Bm8OA
gBd0kntD1Xm5g8KGLk51pskBFV0GGan05sELOMwvfwzkvRcKEq0hjCpFlsmk7gHOKebuUA8EF4qi
h3oQ9VKdlgyZ6jlkYCy/M3/eXdqYqJgq3/3l6ygycXu8K81x2fRQQZel6P/4eLgwT0OcwibAanbm
IyRc+hRJbgLg4Kz/jmP+GyRndT6SjZGm4TlMkyi9PiCSx9hVMKbCei7xDYjWGr45ONoUOW1L+aNi
FHs0t9cjWIhPjQj6kgXpCmQvkmA6v/8PGz+aUXlLRaCjbfxcp60xAMaOdLDA5SiwioxBfBDFwx19
WQIHJWXaieH3sn6dN9fqbby/ce4DOeaAGptlpd+FOMFqOTAFTOE9QHqmMLkKP3QIAPO13cGP7bUa
n8l+8cBo61E7KCFYsJWeQAvN+U865bqECaAxx4ka8I3yjGGnjPKZ57KseiWwMPD4b9v5TZIUxRYG
fMKUCp9cBuU2g6n6KnXUHiH6kgM3GnLh1wmycLKFzPXC2L1cYiHOYQ7lNDi34ILk2t+2V1CtgVBE
w3mpfI1MKis7GgUyRCfDxzPMLuzJ1nIMJtStMa4wx2hdq6q88rEK02DhPxgwNRvMG6h0hW74RZF2
BjjxXQZHuwS8eJ/ylW4oT9B3Vu0bzuqeRLB9jAsiun21dWoYNhI0Eyf110YjISxVsxeCiD7uhMfU
tCN5EEaLBfK3oos9gTs2uBg+R6/rZDXMrMQp+vVBh33sNNrEOFS4dNV5nyH2d0bFgBXsjrPhtzIU
VkI/7fo4eTH1usIgZqvF9gFo1RW+6eEK/Ra3w2pYfjDKADaq4nVCpNUUEE5cTzZ9TmZNUKoZCpAW
7NOr9I4nW1EFttL95ZiJ61OhFEgATylRKaU+cz/s18k1FKtMhflMuq+U01D2MsxT3ORPdnEhlBM2
CU3PchwEsQqlK5a1PZ3lVDgfRdB62ffeWmMUkIc3Jk87p6p5JCpNjCbN+y+ldMxUS1w4JTv+Cctr
oP19nPDMOgOL9eCsDGAGXeoPUrzey4pNV5GkXSFNDSF6I6h050Qp+NugnsX3f8D1EJoloMuZgQSh
GraSmic+qlNr7zKuHKgL9ROcz2cPOrrhRK3nJTw+CfRy9yeKe11FpI4bk2jGbU+nERBNy/E4qrOi
kS9XtE3w04zEtaA3Gnpy/alm9146US+YzbI9zpO0/hEGeYkz7r5i+ayfbzAgRZSqj/fhRf5Fk3rl
OmlAZzxdZXE2mDS13ryJrNRRGGWqS5u/J0VX8Jx2yWBkKpvrMmJs/5/uc/5kgJhtyGHpMwXJ8CfB
/o8FbmhD3Tl+U6tbK/6w5Y9yNZtB9WjjKEGVVXlJsgwJ4jq3C5zuFKCSZu7owznwhDWfQtCcCu1l
sp8NqMFgDnJaNpuhMv0skhtXNYouBPAjEnzRsDXXwmLJ//lML1UABuPZgc4H1JFojuizKXwGznc4
5YGEWpUxt6ox0m7lAyhJLuG9VDfkUieYaBcLSTP1urAleWkxEe9F8Jvakg7jjrxc+D2o6FxfOWt1
801fbmPFNqBcEcBINzQpnvYGRZhfJMaIbEX6DoMVRX6uDNhwRu29f4CcFtGC0hvuzekOBl5F0nDJ
pJHHBC8XzfEXxxKh36JzlFO40O9Ul8e0sYwWRraKLoteS7d6ofVdVYeSVFVKvw7Yv4uN9Jdcf8T0
TJo9NnXLzLlN1Gl203hXvwhlevYYjVoJlBkRWvNBaO1a7SktL3rOeSK9GVTyd3pUjLIreHShzQyu
ctUBlR9ceQCwlom0/qx5pf2oG020Dpp4vvGidXSrcby+/Wjh1zCAJDnujncj3+3lNGRy8ubQWhEY
2frr6KclV/SiECHB+NO5Y3qkkf89Fyz6zaxyR9y1g8yzhwyrtZWuWTgq2CyCsIILd2f7vpVTE1bC
mj/JuoRK/veAcrOlMtfWop4TkInCtlykeB7Urc18q4Y68/Q0wYovX3upxQ0eFW7+XQhcPz5Kr00g
i45YcAxL6qQHVEmXj9dT3iZ7PtGkd4+Qlw7OAR7y6NuypatSKnVGCusmiPwcfZeBuqnA2w4jc+UO
hgds+yJ/u9sdZkE95o1osfKvrceJwO8WKHQkT4gNf+M5u1aO9D+yJDfFWELeksH0yIDjElpWWmdn
U9TraFOTRJLon5hbJmV05Kz/cQhUSjigQKnJv8ZpzDm663TLEv/Xv/TZjNRS3wYqx46EkCZkOVAv
nko397wAdL5MvaTbRwMZqdMprr2aITa4dPYZ7c7n8mRkYIi+1i4x+MCpFrknerc3AW7UaRumeE18
RGXh1hS7mDu5368jftvL7PKqi7tcErHcohdWNlBjT7yr2fF36LOtoZy4eeClrCgriTWZ/w509L7k
igRCIpwiTZJc40TSY6ECjBP/QwjGedNcwL5mqiURuqSj2zLmYd66JyP6zuOTauL0QCEjqKecJ6dA
id44mIBXzAyXItiBBvbjTuGjmf/8wPwz8dZEL+7uoHZUSrMgWsFvcCcZSCK2My7pGdHdawkPpa6l
fZ6GAux+7nSlB0CkeXSNTrkNgw7kcBvoCq5rT4gC6AHrV0ed5O+qxkkiZxuiwfjs1GHD4AoxBYN5
2lHOhlAth7n8cpkjGOnlyzTFpwgeqrtmQih6TnpBktn41LDroLxOQW6+wHQ9298RLlCXuqBXdBZ+
NRooZ9pM+he849ScKkL1D19b/o31wZQfCknRa6nwfOTandBoIe4u91YpMgJ+wCHps/5cBeJ18tI0
LP6C0gGmgp0XOHrMt4NGWuJL97Ddc15SVMeogmMCDrz0n6r+LRNBk2u1QuX6a4HSKKmyp66DiU0k
WIe+NY2pVtdAPSlnzCcZ0Vy7YYjRSBw8SOu8LDBzEGWm5nawCF2Pvv2IkG8IzwNyTtClE0wZrV6F
9kfSgxC3aSIZIC0Cj2tUSExC0TlGvylh5dtZ8Nb7lSek5vgeoFV7+bPniE6hl8e5qprGI+kE55Qu
eFin4gk3yWWoZ40hwxua2V5bJa0niRBNP1WEPbNXZ5TTV0ZL1LDCkJw+CX+OqFJwSLOD7xOdEkwc
MXkCs9LmUSBARsLHZOoK0YExWli7B1gHdq5ZbljtAbNPCcJMknLlcWpwnqtU33/lsskFgN8asQpy
i6reh2uBlBXbH1it2VAIqn314BxKXsRi0ccmsFnnytWibPq5DDmW262sXaDBSyBj/Qa1uG6fUdHj
UVjokpKPhwxwqAQxZp2kGgC7JhTzlFAcNcsdgg7KHWDrn3vkfup5BxdYk5LdxGJh6jehIb/sctYd
ldTcpubEWCjuiOSC0/hFUbaZO/DeAy0qe0ldxFaXaGuDGTzZYayMMGauBlJ633ALt8hpP0PMa8dL
6JosT7C3NHqAKonektzuBV8POfMe8t8SyYeEVyt7gQLZZGWH+zU1kU5Gq/xN4BHt72LMnEZo/XXx
/4vqMFyukfXgKjUHNSmpBpKYwhwC6g1lUYZVxxKpKwMMrN8iJ6BPQ/1dEW12taQDV4RG97tDWR8Y
AaDcp8QOhj00L7lI4ycyfKPv9LNb6AbpBt6T8Ohlhc827zwXAVbpc5WrdJQGz8TeSwxwCc/X7a5g
qd9K/Sym90YgKi0H51OFEydSpLx5EtdRtcr8MkRtsATS2bzh5bhguq2F7IkfqdLfyAZ1/YUwJdpK
lgykY/UDXFrqvqJMLCPGP/ed3LCKbgPf3SoNW9n1wWH8nJdgFoH2G0TFPD9hTff3bpIEeqxvNLc0
o+Cv549YzMduXutPCXiLWoz6VQE7oktrkmm6SJfVGgrJTtfSH1pnLONSYZz60SbdG25dAD7Ix3wy
l8zHiUSyHL69zszk8HBluPrj3j7mZJLEprYEEG0pGqbBq9jSiyto4DRIwMYbdY2cNs3BRhxDlHPg
2k6W35D4iQVe+oSc5mDoR44AeVq5bLKK7aiwWPxeJ32akIg8Db5wA59Twe05GXGjKqJCIC79Y92V
Mlj9GcTs3bbPkyKSkIeO+cfdfG3KPe+EpNSCJ1AgJ62r/Dl2ikfUDsOaBpK8sHnsEV3m3vyX1Zwb
BA9n/Lx7o8kty36Qjl+Xw3Azuxd/hPRq4+2DYOJT4mWKdyGiJ7ZfbWunY1NVAnOuzX725LcAOUOw
BBF/i2qRKUi9xp+l+KqTCPL2tU9sGPThf+pOPOeFgA825NScnvCpKjXtEFFWOSlH+nOZfMC4NAgy
o8k9gwE34paRB8r8eZ/VrGH8sEgApmpUEbWRjOCJpNI+sLABnvABYAgOyf9XEwEjr4geYls+xHKd
uXw1TOYMv7zEnZsY6IVZPUQ1wQcl1dDBdcQK8Le7RYsLi3xmlnLzHd1CbHG2o0KkBnouUefNm+ZX
rQTFtz192yycrj9t4BdFEzbkjChhAFJWNDJ6qWQbAoRFULv2WTtPa7t9DN0WijpVJWG3XslOBmdi
KMrxL+RTyLjmdVugS7EwhRHzigAgPnaompiGyDQvYZoRbP3GYSHicw7CnVeOBgSNth+QuDGqPP/l
LlJkaP0yIIU8ZQOYtMUD4605wioL3szU/9+XWwT/2+kB3oxYMVG7couMKx1BusgCI7Oj2NJHO5BJ
r+aIP9vPrDdlatieuGUb8/BPgopazPJXGfBeW2eunw1B4kTd+IoasSYENPqTUSPn4R7zpeyNVEEF
fCDZVjBMdI5TYLVTGF5+nzyezkA3PCDTGZic8iKqubaDWdTUvAFrpE7DBnO63XUyChZGLG2tq43Y
qs7KxC+yy/ZLqqy9+qgfjjHm9qXEB/jtQeSkcVoz8flyxl/E8MvEJQ+nPkakOa9D/L8k6i0Sgzam
ybA3Ybu+1VN5CKcFdViw6HCxbl1U9cArYX04CLWaf2w+0XfLq2fiMw3e7jErZsuyXHG3LRw5U0sW
3WnBngQfKBOvDnIqUo7Ggh+0wxe6VPEkPLt081BpMU11DCJ5Qs4I6mTRGg0qjeJllyelt01I52TR
1hANP9Aw3m1NVntxIPpwzfraghYDyIDVlhAClsaFahUpo8NxS9H1Ex9m8/BOqCyoE3wkkz9jfafb
l3vN6EjtlwN6UXIMlPU1h+0pMkScJoasL+kdb5fLZwkeHQCFXreUjIOzW2PwQ427FcrSwMWpbAB7
9bdsPI2tPcjfVo5MauXyUrc2YiwujDDinprZmWxih1bSKkVhlesQRROZJWd5/ECZ0UKtxzVwp2bX
yWdCy0Rx+ihw/QikMg4uOjcoeTxzG+biTt32uSQCSM/fypWjkS3WdzeAtFl91EYpSQ/sVZFXzmmQ
dkMV5ASpPEQ7ujRJTDJGygqhmVj0AKPo1aqlUOXsTH+UnrIzAwhqPZMNm7YDIklhTixSevJspMFx
NgHFNmWBuWw79lrUVdURoBQwFo1uL67hk9iYZxbcZeZyw9P4WqwUYMPZBM+UVuLSZcPSrZ+sjOoM
mV+hMmQwBuANeK4CGbefYhzFT2PAfKeL7GKFMllADRuwZjVg7lM3fByiGzaAO9QNlJIfmuNBQO70
ylxk4n72rHCiE0WgNfVAd56fEDokBi/gfn+Lj8ancZt6czVM1QQEGSi/JC5j1u5K1xHVvqK6XbhK
3d+rmMzLUkS31Pv/txaaqUDFr1EHtRnxAmiMnGu14hXudeG+dqcgg3E2eEWArfFO2aDa9J4RhtJx
cc9Xe49uO4K4CDeiMrzgDyH6jp95TpHTTGsq4JwxzVuPp50ELL+zOI/ZKcXckiLeM6pP30NsSjq0
Uw5puKXUBOylbXtCVmqKI71zDIgPhajrrbqrxhIQNPc1XaTIFLlgZh8BRrxgtXc3dOuJ/KhdmQ6u
1nSz1OuQHgivyYLvxTtWUP8p+6kq/cAujDAMRABVe+99UN8td4DfhoiqKKjhBsw0BnXptb00u8Lq
TvRByv2sZs32E0t36cUHNrCAkiQXiGDl+35lNoHnM0NVP7vx06rxx6LCKsyCORJmnQJNeDNpn7qv
K1MmrKwGKDWi92P8EuTq1ugibLidrnd335Q0TYK9kHUBSbPYfn++4X6XIrogLFwsaeZWuRYS46jw
ujE9AUEpTki9yImBj0PnB/6BHfRpSM3UZJOax3nI45q+g8xaK2y79DAHCDvqLpftNJdZ0tzI4sn2
L3S1XdXIGLlLxZ1O8nllIJBd3UP5BsRSHZzzIw5uM6F3KYNaZ0ECGgA08M5Zj9YA0zAakFgpMn51
swXf9xr0G6Yg5IqVEdUqydHQBUtLRI8yNXsZEecsnIfdMiZuEWF6XDjMnPGlzJMjWfDt6xNG6OoC
EctjYZXrOlISVyUUG2i7c+WW4mm535UrM2eXdNtNKoVs4UJ0/OndJSUNpFMaOnlBOPsNj+q76iGz
r6njQZXAuZ7/jsLMOqgnBTe9mUj6HtkNkylZBPQCVDr/zR0bGF1mxWrc7ITElZ4zHF5tQT6ClTSW
qeuMryEXURG5CA7n9EAre4JecWnnbC0kpKEz5x7bLl6OpsO3kr91agyBVJRX0gg/I6r2og3L7Dz9
6sI6AMbiGKBriHfkJWzzykuhMrjmZf09wM680hm6cdHvmL2JUs475yLPvniZY1Bu/q+Iy1V6bM10
1uapFa5v6TJgtfns5B3Iu7hB7EqChBQeDm1I33c5I5O9DJ/V2IS//shlVognaOvkOUonfBbqni/W
kWhPLRDev9vUUYY5W1ZjgQrKcl9+Ss3Io/d5W9P6YA9q98idCUsUBzaAC7sklsHPRo+iMGoYfl5c
Jn/o5JF23GiokPoLHBLV98JeVLAhi9zex5E6HgB/upmXjgza+I4s5g1BZwjt2YHkLSyJUTpiHKoK
zF3whsdySILqMKYgvPQtWxzrI/ZP+cRefCXlITyWGN/PJWsfdEVKxveLNjSQf2HIoVBs3upoDecl
BNuDnfTRr4XeA1n/rN+8hrFUFn/ZA0g352sUnfcm80TJDMihfDZu2UGlI12p8vky9x7gxX6pLg2+
BfszqY2UX9+2do0S0OX0czVr3fi9NR21c0te14otQbkeXq258qa3kjmL8nDp8SwKFAE61yo+39Rl
aFQcit2iBhGmlKEg1O1mjE6jG05x+II75GLKJASehizWMLECcojY9gT0jRDCoLKjjKGX3XY9VYgS
fxImNPIT3yDryE+LWISk0KVmtwkj/S2xzSIZXHWUzayUBRZi1K5eTj+YifaT5QJc8buUxZt11z4l
tR8mO+KhYbAl19OyeWanbWCdBazt/p/OYBhH8pY91qilFZvRctXLEA8LF+6YcwLbpnIwzYwEBfDv
4PTmt1nC5pjJN7pAoar/bSP2c0hYmjWzYGnxrKzHCiFPODBttxJy6+eUFafv2BvSdpI2UkDNN+tT
bninNxw6/9ePKUoX09SlzNa9NWlq49vyxs6MNEvw9oqeFY3ffgsZmzec//PkeovWASTwfiJUTPyu
N0AWxv+PX81C6F1QzGjaJsblTu6G/XWejj+0VZmAM666/f3NspzCGEUjGHz/rijz2q5k99KLRLhk
Pct6BxrzwiIMq0vSEzBRZea2peqIMXBV1xbq3MdrkLyGsn7dokM5J4ymNR1reX+TZtgf8P5HPf4m
2+UwStOgYLDBbhwH71U9RMqxa5jGRLswPTNLmbN7TChmd5zqkvPHcYjnvnWEwu4mLAPeYiEaYapx
1js968ViMxO5/rA2HZRDBRZ47yw5Ymzwz2WgNTASQ39vJ2bqqdFdN97/pQNkccvUP51B1d79IAQX
OdkOATHNa20KDw7rc0OYR09pAdu5klS5d+htOJdwSNph06gDoULkXN+XH80GJipyH3udP3aqRBvP
CDBHeCA/dAdPJqSXrzvm5qzVBdaNcZ0b565Yn8WjiM8CJ2nuw2bP5p0bRS4DnG1xYQlEHiDqxb1P
PbGYn5/XS4wVabaBZ6rRRjiH5I4qkLFVUm9tGFVCcbVPMjUVF52V39KWUez32M+D50omxYgMSIBd
FWhL2Y7uMK1D8fcpg6fqgYfF9cZQmfEPJFbRcR1eAZOW3Er5pF4NAxarlT2YkDql26UbYRfa5iFn
Bzo27QR6JUzQgiesK0Guqf2YqCfp//FZILpXwMGScl8/Egaj1LxhbPqlaMTgmbajkTnvY26WEI+H
HnoPxB21Qz6k52QKLCh/DGFZlVFktsLuVclrz61NGhjyhJIEvYSZ4YBJ3NIIQL4z1chq75jYZ22m
koAgBZyckARM9JfyrcZ3qEJI7H9mswZwNYKgRZv5254R23j8EMyw+sNhzG7EeFBpslrajmtyhcBl
UJO1UuRSPIRCQVC4NijSZVxUm4CcWRSWn+Qp4b4vbSoipC7xeezqSt6qot/JNj5YwF1iwYl64wLg
55w1Lp8wBAxDo2xytiF1pzYsumwZtAsXXpKM0xbINO18c/jZ1pqyuZVndV16p3goBeDsvAmO8/LA
S4VsLBBfwPJ7K4/2wrpJwWGfVjwCkiRpvAKf68TElEOsdOolDHwU+jtgitPN7AlxT9tuw06txy9a
tn/B+GneHG0Rba7DDHotqlcxXr9P2qXGyOZkubMb0LBXYiFZyYJciR67JBcTZQIs02+OEeK7bg0b
Y+EEHtOeIK4X7tYCbeyBtbTH97h9uU6nVbhoogYedqoorn3SFUU5TJz5MQL2niojSag9susH2Onb
i5f0pXHNXhIQYhDkOzkDZfnGFGYa/sx1DM/yLgXYo1Bdh6viYUI/YS2kHWjeQr8fkuDlg+UKdr98
GU66k7idp9M3Fz3Qg3TqGdwoDSnxuTfJHb6P7RekQPnwWODD628Nj5psLCYRaFQIqvXO8H2WTNcI
6+tvFCiSjHv2G4zMoQaBElO6b3X4x1GrVfUDsPoeiFDgavyAPmBD9WzJdyqnPZC2mBVRKnOHS8Sy
HI8JTep76zMtP1lbJLOX8dlknO4G4gflr8+6yiUFTVdd4SlSTDLeqhHjaAb1gcIqqdGlRyLQhywZ
Z78JdcbxUF3ovr+4Pso1ImQhJyxQ2v1KI4C1cPoawf9ydjciD++XnMVkQGnF/6pLscgIkd4Pa6Xm
LR36C2XG3/tQOFVk6Wog1mVjYVWGkMYnzyRgJeUlIndsWeuC7RrD326anlYP6ml20YdEToKlsUTE
eiZRgoz2WM+1aXb/0MlMFXj6m0mWZvAlhXnrPbU60qRI5xEESpUv+tMjs+cOoUPfVXfq21VL2aB0
O/fkjH4LanZUthRYwXvANkwCtH9buRcYCZceVeWVgPegp/z1QeejOJNS3xytQ0L5pic68/Isigo3
PGQGjxn3qBemp3KwVqIjV8MnkjLfkHC6SFSdo/0BFaSZ09YaPF/AF2SsPUP6G9iv+BKZbxRatuqT
o85tAhL17DByYw6pzDEd3A1wKcgfu4lY9VAjz8YM7m52jNJ+6GyNP7nIhv5Qj8eCeoFUbpPyU3vY
CVkKcJzcfoCv6E9LfxX+Gx+sB0/j3DvXUTY/e1iYFFOvw/0ORdQmX8ZfdDBNt+bj+NWuahg4wLvI
rI8ZJmUh3+/EheeYsCG08Ijau7nDBtjAotx+M13mSgQLdxkCoVmZ7YE5sWkr3SGE/8WG1xcbCtrl
aZNo5aOumVfoFkwopemUPSX7oS9czdXVPmAhHQOLln37Mnbl/KFcbmNl/1gkm0M6ZwfPR5B236LN
IfDY4hLGC+hu4Y3AbKFHHKc0ucoID2FhOhbAFTFySDGs5gaZGgjurCSZX13Mjz2NoN64ph7AgJJs
qBGc+3xd4bKH41BGf7HKMHeB0ALLpHv8n/HqSE5IJ3oNX0Z4eFXbo4/xCMM2tob3l5aqB/sTTGXg
0ziYDckp4JIpnIw2fA9mJ9R8BY9DYmlrwcGn/clehU6zwBYEk/hzd5owX9sghE0Dm9BT0RvGpcVL
ycH/xt4Z+xi4unL5W9pGHHjAZ33l8jk1qIIWZNhZskcRTtBH3xIWH5Mt37Yol+15Bo35A/dlU5G3
RuFUT1TEpT3DZfUj2kkEdQzbDneIWLi7g0cFrRJuUnPGa0sBLakWLCbgxm1uYErIOQXEdhrlauk6
7SSvTtUzyFz3/qySyYVbBffmyoYRQHajYGa16/9yMmcwBglsFCH93H5J8BoOPnUewjmRpwjLI1h6
7dHLB93RwjCy9B3pRfXvUvK8ehwiZuHHsAEMT97Nfh2lY9bf08yuaFx4mWCE8MdgV1xGeWBJ3Ckj
nUvyD0an7oZIg4KN7OU6adic76pIdcqFY0tmzdNuRc8kTR9yYdnN+8cEn1gnVptki4mBFearoxAU
boYVg8YqyxsqWRXz/AK3VGCPOyLF966YxIRKD+9N8BRPRj8ov27mgNfRH4bk9baHD3gbS43up7oY
4snFh2/aJr86qQ87E6qpYuI3dXc/NjNqN8nbrjU7ExkJOx7CLq3sJ9b4J5HUYsp2Q2G3ZmD1BQWm
ikn6vvF24UksSLhOSmuiJS55ESHap0it3I4DmR2f94O52fX1zfS2UlmfXBqEJtqYmZdqAZuGNZ+U
J9KTY1FEF//IGHpSMyyNmFfRj0rApPZT6sEEySkGrdLxT4M1rMufCROsxme6Be1V+v2efQuKs/mK
PxuctuLIbx3duhnNr8CvuzgqoQY1xXS+segsSeiBQUy0kY0W9/Gh5lMgEPNKSfToEKCHLEL0cm6X
m+2W2Glzm+kS+tBEMFCVW6aEcNI+8S13khpBFkMIsO6TEba/tU3IO8mufrWEcxAG8ZBW9nlfUwMz
CMWraG4V2ftByk286VLoU3DgcuSZRkwZ+nOCtCVRlpXT2D07mz6OM+Op5+OerQ3EqHzYEdmsgzbL
ttA+P5ZmiM/uPz+gRJHUcqeONDhfzEhhkqROkisH+A401cbB6d5E70Z1IcpyZDKHsYO4UAotDNBC
hvQnylDuGWoOZ+H7JOomIsInTeKXdQ1+QLhi+BLi8tookwIKM/CAHSiv1lLl75ODUxaXGrFBTtbu
j84quZOzS0rmIacgz4KdAtHwjr+zf+zB4dT7oUgQWfsaniLMQs/8F6A02+fo4FRt4OkZ7zLnSPlH
HUBLVyAZU464lqMcsgoWjQJ6A4/uam2jG13jgNQD/aDzc1sYGO7CLkR6dYw4hxqailXKCHKfKlzp
IDXKPJh8GTarB8/e1IVd7DjpdIkISQOv0EFTrvt2V1DH7XsAyxbq0z2e+75JvRc5La0g8/rE5PyJ
VFWnY0FRdBi7Xe5NkNBk4UwZpmKMHJLQl/BD092lRtS7FuFxKgYwEN2N87WJBagVe4Pkri60Ynel
UyXeyiWw34xXoIaX8BI10tO2GAZO+EUZaoV1pe8IaF8zGr4d8iQ+ObfAVj+pCS6NySS1CtyLJTpE
ajA2cgmYoHASTbshNncJbdEOlhIXnwnUiru+UVfib3bBtWUsPL5fHOP3a3lsrDpt76+ehrnnk/bd
s6yR/zk0HIrj9NjmYVU089S/x22EWka4LHcaK4ICODQa7FDPWSd7CKtYpkOjnceo0EoQN4ZWGvho
JsYQsR0LzG8F3BOwjJk3UplZUmUwamcUeOTTBzQULOSzvIBDHDpWm/yxlZO9SHVg2G/aIeuEJW7+
dPV3BG8ITiSQTXLQSr8kvHOG59GIoH+aOrydayZ8+nb2EDW6faZ/xuIyT+kdRgWNPZNFrhdCQF0E
jwtCWMWZJoCO7Dt4P3ATsPhX3t0uWKjTOnkPZWOMIOVPPLRJYqlrpm/XGgA+u3zPO29DbZy5A9Fn
UcBEi4/P6N6/0ZNP3p52W8Z768UOaE1t3c3i05Q6qMMRo5J8GR0hsjlZDx6wIKDDO+bOjarQX9T6
pFTl4UFZx/g7D7rnWcBXU2Cx6YzK8d4G3cLbcec5Wkup/Fq/wMbfeWT+aOKXn9CulFkun3EeO2ZQ
jCkFs68lqiwJvuqBDyYDb28+jPtVkI7vq6SKFJpCSVOgtJiJ5flTW4YkuXnGVM5tz8OSjZZL8xIm
y75F7BcQFPu7+uoJE3MlPoO5jjCph5Ym0KpEq1V1a3lbAvgWN+VqaU5+nZTUsg5K2RXiwHz2dDFY
UYJKWDEXcGPUJHUVVA8mwAwCRzKTFSBqqcls7tTKC1zHgSyKEoxpQ6IttqEKOVQ7S73+jkgwPNj9
KnFRYJLBJAw6AwQ9ZPY8D6hPo6e3VWHXHEHOTlN1EmPSDF72gF3GqpYRacK2uzMCi6d7dv/NOs8w
ji597w8WEHNdo3YlUYEKfzHpZURjNcD4WirNKP+hUeoMgayaLg2VKuBX32TrSfrjYD5QJUZMm+lW
9QEMtOPPJTz97iAgtlcTLp7ZOuCOZTjnjUavmHOg4/FDar6MAWMBGDuJ+NRe3c9AD1/bWn9l9eLL
7orXX9fmVePesk6cP5/qc8z2GDTgidpwtouLdwV90vXLMRgZA8ulzcWHviUxBy8Ne9bQQ/lZdr8p
O4C8epaDRmSg2tBpQYM807yolvg/AgsWFW95rgzGqDA0H8pfv5xvvmD1dChvbUgfJjnRtqsL2Q22
3RgxZtGZtPc3HjpCpzDTJ8fxCqd28hVtVMsR1DAl/DoWc9u7ORgU13mINSM8z/S7hHvFmgdpUqKV
zTs0w9Y7iiEAlQJTePYapVhpABhR7cEfiPle4qBExCTyNhT8jdljTmp2lwQ1DQSLkP1wz5MsM/M+
i70AmD5EtOuKKUmDJxkE8eprT3FxqsyiAjTuX+c5y3MesBFbcE2pSNHFmAKsntAv55eWtUysy1yu
Dmf+owIVe2sfPR8AvfIiVeYi+27Ibu0QS6ngNOG/wZbGOwnIo5bbqR2vGuCZ2SW32EPqL4XzUU7y
nTiBZ7fmSFPpUFZBmpuvOOBhGuNRT4A+MGgudD8QHujoMJXUaDt2dDPrkqRxi90O8EsrqC8mjj0k
1cQ8lXmC7Wr6+Lx+99VCuurnC3sPQUlY6Y2O7fS9D6epQuPgSNkgJKyH+Zp0zoFA7S1cee1CqOtZ
BhS5VjKuLVRclsqIEK+y1qAk4EknoV1eKk+8hr6R0yQ41UstOsVvc4KZ7YMVCF7nIC3ero0ULb30
WC99yQU9VeRza4roo4atzSxUglLgWDI27FbcFE3Yq+SmR2M7NYkzlbNXnW9YleYSxMyGXbaefrif
UCwLXjbiJ/Kiy6LIc9FzbZvicDSbA9Ph5nfr0MXIuQQlL6oNxr3HAQO+e65ye7qBpnFm3CpryIAD
PajJqsiPk+qBxUwcMP6LXAlNyenfU4v+1/e+SbEGhWB9ZHSbc1SRNWyPyDosKIZwIx9vXj21zDcs
mum88VKZkXF8Y+zT5fzTbKgUdicpFHW3x/11IN2m8a8K3kKmoQ/0Qa5iUEF7LJGY+8alDQlBfCFH
uJOvJId298VEnV7YEOaUEAqJmTt+N3jQMgNd76x0/RgqmFTuxsQcCFTDFc1RfBw4PbOQgl5vOKFL
MvbagDtdAVxbhrXOt5DmqW0mPwFd5nYZBEfXvuaaSphzMxAJnqhj2xDzpr0w/fXIzUnXujMsozpp
cbQML5XFx20ppMn3WO5098eUEfXI9YvGJQZRwU8kpjFEmB/gXGkZmM/7az45O5mQ0jAb0RazH4vW
OKR0WbSSSSeXA4JbuvQArinni4H4b2CFcQvI7f5bem4zORJf9QcVjpjtsxN2HxE3Xe/deG9BEGG/
lVUgJVM+nj40QJpKeklhIqQebQ23nkqXgGP6MlD8Jh3kEfZtUtDu3lLm6rW4Rgz44/1AP1+fxTtH
2qFemijQlk5Gf47+2ZeRrTdAfQ4BGcqMWydgCHsmMLSMql5GWr51yobHkBFbe57MaC2vHMDivo/4
vDqkmLv1IK530YC8tMAkyRsHILfqOPYCLkM34Zcj+uPdDztnxGgFDONHXsO0Khd3Hpu/laZGDpk1
NvEwX/flandkcbD4LnM5/jPos/l4llxtIkjHeOWEGWibksHXC+Y3ztv7BpOX0usN3qRZY8suh7+7
EW0HQapnDh4Df4YAVwdvXKttuXt7YxMo4kPzjf3Bo9QSiBwh7ovMJ1IqALR8nCMZFEti0aqGbOaO
KUdh4KKIAHjN0newbGOnyLT/1C/PKIcbM+Fa5d9sCDkJ//tf75Dc09DS4IagwYPJg4YZkxlIsOFG
ghYWdRo8Ru0Slfiq5w0bsDaOFWqh8qXpisO9ARjt0RzQUPQ/bxvDoBHHzA0DYEChGQi/cjzylASo
ADlBT2MCVCQSCjAZZvofTJJrUBGnuQfDWR6C5pCmRO763NnJRJzC3HGsc6yBE6PwjuR5wyFN57UJ
ctSJSauLFyjWQcciSWc9kUjjt+PybI9y6A9rADOk3beH9OQ1R2qZvfbCNFBS6vdVQ48DzbJgdVMS
kIXcP8jxTILIb8kGsJi+zlhCH/bykViZ48QLYGV4jZ7OnUv4MsCi2WvYFMwApreEesh21qLriVg1
fQ0zP5Si25SqX4GdaTIgEIjSpuUkcNHdvKeJ30XRup8Bo/qJLLDu4GR6GLU6eFUR9/V0SNklnPpw
xA2uNHZ2DD/S64D7AAMGmgmUm5r3hW0pxoGafrd67QDqRFhvBC4yuRu/KbMjFxb9oLjOTQSv/7Hu
TZlyUOsxBO6hmbdmuJap838x7/yG9K3IP/xjuUAxAZbfCckcBNQBPqsZc8aSgdu9wV4VyjUlXncP
aGQ8m4Tnh/PkKH10cBldpcGp/brpS98RJnt8hrOLTLMDO60aLvYwIm5tQ2EW3ct5l43Ks4yB0DGO
Ohvi4J9pftS5tqY9ds9gu+Ay0rNFUnwcjlVY1pcT7F49pT+9bxFBGMfcpZJzSMFtSIc3R6h8EV9E
2v5fQlPIxQej02pQUWkpguQThY7Wr5W7yR2JGH3z8cuOiS0cNdkJ2WMnb+LL7cZP2N6lPLh4FrSH
m4kLKoYAI3jg7viEj/IitS7IXmtQ4Gr9vRHA53oBVrlpcE6zTZxIYTMaqaVPZSwKvkQl7EVXno51
S+ujzh2W8dzNSw6/RgQ6SpA9mt7mgsWCuNyiaO5pfHPFO0LgHB6bjyYDb2CZ0MdIwJCXyW4Ekk9k
1Jf1m4Mj+O0NhU2Qd9LZgJoNzkdmXEGBFFZCslKE1Z9MzdIT3+Mm2Jg4KdWBJhvHfU1jRIWLZYHg
sJ9RM/0PBxGi9HadRWsX7ALQO4r3Mdrkyc9uvay3m6kviHOGIu8wBaprG4aLGxnMjL0XYHRUM5N1
qdhGjXjHmbs3HoVuwJN4thD6w5uv5c3qMhXHBSlsbQeeANYASQ2igo7AhZEAbcIlq4hXJEcjNn06
idXOQaRw3P144l7mO0LM5mR7kcuOC8t3oG4F1h5ALbd8T4XyTECpL/tOcoyXVTj8DP7gikRX3vJ+
3R5zxHIglU7RYpPWvrSDH9J2NbGwX869KeVyLjsu2mb7JlTljfrIphhAmWVofYEnJ4hNfNCCosWC
30M0hqcULN+5ERv32u51f2a9qsdcRRYXemzdHrY60mBoLFDTZTNkagb+TcTizLdLnFraM+A/ucZO
SWIX8UmFubdy+VIJsqsT2TOEz/nUIJdDObAJCQVVzFHTWX2Nwdu4zl43u62vFmQqgjOreis+n8d4
oy2U5nN8mshVG5Ff0yIw1h2ILoIoW5hOFs0SV9OaHhq1Z0TUMxCVNAeYQ4g4ZBYiSH9WIHq6Nh0d
y1xqg3OUGam7LRstVsj77KqVo7qoUkC/iJ7u7uz1cYe0/h8NnnUPslfCY3ohTLVLwZR6/feiAGEn
Ghi83ZJZ0Eku5qfT8tH/Lk8FnFlqiRXm7S3yfX28gAEFHPRlXjrSZvv3wsa3Xpr8ot5xq6P9ymis
encaWwPAarqpWQe0fiwCnpBJvhF2iw6b0aymH58uCor/HjonrMuRUpRkCKdTBglu773+SC4jghVK
bUayLZrETAR8DkS3lDbYwCHGkgdw+JY9i8VN82ObSC8tRuO22Pi9FETOFsmZ8h6F2eK2gV9cNH9S
hxE2CqYVDVgLs7xQs8VdB+djSe8dj52JKg0Qa3fjVZcOInXFq0IdIrs1C2Oyuib+Uxv0m/YCqoH4
slpgpbZ89qKD0c/eNdVYyQJKNUOqL+Moawxlli8ABPdBXIg23eeL2nrdQ7JW19V9q+C+fSpqFbxG
2Zacth4ht3FB5OgEhKbOEFmy34q/cihCNbwuAF7FODCSRyuP1iUBOpMWf9DzrWyFAdxS8vGt5C7N
mMjMncEdL6tIAKzINiXYL9BXXLqocDrT2cPjViHYPI+C188rxnhQXwAWG/nVnezXoxVsm6ZD8jS4
6t04XaNMk2ku6zdzSeLPodnsLxXXxE5Bz5VtRjKZgO+bPEIjffWk+0fgpwQOarR8nmVobFkfXYlh
BRcaPgoDTeANEbgoVslaJagBTaMWrzI0dErRBD1py5H3W84Gc9q/80A+m7OD+Ot8riBy8vWrc60s
QEeRZoCXwJZYLbu+yQR2x+nImq0l72wjsh+RFgZ7gfHCNcvf3uBXgAfi7U6pnxUWFeiRPWobqHOd
qo29lvE4cnIS02iCQAyPimt1EzBfltCNnnPOd4A0TJBIDO4tU1BlH2711Az0hiwfvlnMSYzKWAJQ
LRzGBDyl+MWr+AL+JsK40k3ZEni9oH1jfprMcwK/ZRiwWYL+1IXQMuvt8OquOS/gvAObyjmj4BVt
3Ufnl0eGCyUp6RrP/Dr70dsdJOnSVOXKfBBoDiEXgPOjxDRg7sfXuxNDQbCg28tG3e+K/sQQLMce
hDbUEdfNA/RxiiVH3JAEkIaRx+9HGZLkk+BjXeqyFTQQIv6HBlGNJhdguQK6q/ppj/YhaB1u2SiH
A/2HMXwouBMuPInyokZFKexn3jpln20aze/ZOuPusJLlyjOUihAv5SLx3+aT81WNfjnjVLGD+8/d
r1DKv4plrwISNneY7K+dfXeZlkC2B1Hdi5NwBt07PT48KI1vyBVtD0GA/Ro9nF2dRQbRRMZsqQ+Y
OJxns1+Ees54ATXZcuAGjIS4kAz5Vjd01DKErMBmd4TpWiC4kcOZSrhSJaaFs3zaMYbL45Kenjgq
ImLM9hbwLfmZBsevCSvkOehhw6D+E1clk8i+0JsdjWqj0DTBNXhu5i9IXT2ajgDuNESyvNlquuJ5
kUyoyNK7E1L46qOjKtCMD8sXLPBKJYmq2OoSUZ30xKAgMykh3U8fYArO0qdysJTI8/zKlJP6/vHO
QJOmgM51UlSNkFnvOS2/yO11QVRqumL5xH3F3xygpFwwuva8JeP3AGRrrg4L1DH/Fu4riAbgfsw/
RyG0QhMge+bcRBbtK5Vq3AjyZn/u3ym0AFqnbWnZ+gLuXiIbh0xHL4x3xiYw6btvbm/xC+Vj6c5Z
dLFtN+pLOtjY6Lg/ltdKH0MzwjUjEBlR0nCIxIPA7MVHeMdwtmO4gfNiAibIyTmkr/Uw1whVhr5V
iqpKvCKInWrMlRSTgBFn6/OKXFqK7DpQtgTEl9OcdQTZhN81aEUjh5Py+FNadboKV3WUW3+SoJiM
RWDL08pZFkadeKMFCAP1SQ+EEdaaRJ9q1cOG+MZ/8Txu7Wk9V0K5zQQ0H/5eHjp79LbR/D5DYtEO
l4fKuUQjdNvngZbw/AtHAVS9Twz51VhVgZs13FWwAk1gJjj0QgSDp9T/Kbxcdhkk434kljEZ2hF4
pqlOGnhaJ4q/JlrVaVWxIHjSndcbyHqcrEzLqmVLtebfflCAUa9B4ssXLi2HTc1zQn9+dqrG+3A7
b02++fKcrqFqNt53PbnOloJQOIb9NuDEeB9RltKHn9GMVS9v0XWkvar8iR7q7zg1D8EMMhZx25yc
DDUzdDplMiF1osHCw6qH+loBdiWF8RnYFx2BWIRaqWvyyJCFnvcN4LVsoyDrjCpv3IlhkNGi45E3
RpvcKvCTLnwTztvtmrKR5eX92FPslsKFuZe7G7RmCvxApf7P7sLXP3BkBcsDzVlpTe6s8W6OFa5I
45hSsPUeEIKrI5Z0jdmBDnlojk6Vyu4YaCGdy/9xyjPKuSz0UU6+4Eutkuyr6TRYDufuLsrpojK9
Mn8MWL5eUGoHOdumMHOwbtO2JRn88lutvg9dju4KB9+58GbDDMgD6xFuHAjn2z71/C0W9RR6gk+V
ePLHRbSshVQ1nDheu7r+aBDpJJiJmwk2xoTRcwSnvGDAaHiEWfpLYb5CztSlGgFF8/LSglEts81w
NKeepzHJ3LKh938A6kvjMhJHxfRorfqfTnl3D8EuWOErM5AtgypFB8gCAaIuHEJsJsF+sMYvT6n0
IOeTHKgf+X8IJD4SKVS8LF06S5wIyBBhvOIy4Z+keygEjcjeXJMdls85Nz2X+Rjksy7ru8lEc8RW
3o1PVD2IwsrJYjzTiuFiYblhRr5MPEhrZQvV//QZE/36mZkS0PoVLwYXt4lao+yIaeSDiJrMyXwA
STbgx5JdL7/aK5YjnS+Cad7PJ1d1It4rZkMhxHLswJSQPoGExDNDquDaehg4cEKuZgM/IcdUCFjX
0oJbT7ElMV6Ddg/KKsGsDgH3/ri0R6eggNbZxs6ThPcCgdzny319VoOBNx1AD2LP5KvSJ3PBZPxM
tHMPJVOh71HebkaxL41kC3SOLrBYl1nMZ0RTBUaAisrIoZ3blxem1uI3nJXQkwFpBeDkjYjljmgU
7HXrIaw1UpBLnzjMhcYiYzLyrztTKFQBFVT6D6pg4qonxbpgQqAE1ULgdmYtYIAt429MpllyZgJW
cRCqVq3cDeyqVayPIJLyY6JFdt3RqvCyF2BoWYq9mwwgmFATCsIi9amWVFzC/WrtKC3F5wPDoJe7
nwIeU3aEB9aLw0GUcAU7gtO+s/+kuG6q1DlpqifkCrREhXWIGs9NAe7cQiJoHn8gcd6Me/mm4MDp
bEW1Xjytp8XJ5+3LqvgCzYUTD/8a/xKE2kIHkrbnqye4rWkQOrqUKgr7Wr1d9//HdFhMyouwzlOw
oviA1/qWhzVLIdwHh2MtsJfGUJzmUbQ7m2TCNce559mls8khvmAX1aZ8wWs8UvmiCJAq7Rxn76Mv
bkLqwMfD4As+nYmnY9bFVRNvnzVETLhJ0v2eMEzRSK2nVtUEskCA0+xDn6uoc7Ln+2WnD14eAaub
GsJOeZqCJs8whKkCbnbfTgmMdz97C5QFRDoxnsXwlXaniHQSBoZnL8mTx9hGDsLOTWPxuXFkLgew
xt7G/sxTVB3XAtfD18lAKBP0Q0FgYRlBrixpvmjoGpqYsQCuRRj2KPOSREh2Q6Eg/F5rzyW3wcVS
ZgnNeM9s7QMQ4cdKv6QC/7um94CFCghdCVs/YYkIpyk59pTMu9Ol8Yb9spCxLuHPwAU65RrHAjZW
r/IIetBFYSMoI/NgmWkHJSGAnI9NYI22lmRMBrp1jaYEtS1BAth6H/k7IfdTIQ2pbIFGBCr65lNl
I+SOKc0g/nLu9NWhzUWsP9gjwyzRKx7UkWcXzsYgkrDJw/gi5nfJAaSzB9gKaPltkr152NvYw0Uv
RCz0qO8gE19ckuidyxMAZTAWqIis305iQsGetocvTU8LXtTcy6qxIjuNkKCLNv4hyjC+4pydUUVv
iX2hbYnb/LK5smNR3l7CM5Rxzmt8kZBUvw+naB+V5ShYFBY/BT6teAljMSYvgbut+h4A1pZxMvUr
RcSKfh8mdfYwkIm1gG+Cm/OBnP8ClHuKjBvFs+PenIVkQB0eQyDwQ2MGIcFcHFdme5KlNxybKy/1
4v+CcSya8D2THKYqmwUFF1r9soMTH3Egro79Yh5KxiCKEDfTgkDYpXVTlgnYYMdJvooXnRIb0YYC
T0fxyBIKD1nGV1IH0B2R2Nm4zYMOsEOQZo6Gugcv7puYQ/v7zQ7Qltvqyw7QN5ReKTelVaTQ/GKb
aBuz641ppWlX3GJgDrQWrxwKn3j13A24k+OO2FprSaYKWntGbPwzAtG5GeFgFIcVbGlmChLL9CtJ
+St64E4PGmZsjr4z6vtkmvqTh9QMXsMz/dDwgL4INV9wXp6oDf25mS45Zbz2CmTUY9vtHAXLmFTn
QSvVo9u3XgDfcLT4UShabQhrYqKNvvQoFZVIiFWpUAbSa4AW/f2l0kI3bpgOxUSIQsI58GLLSIR7
ffiXEsNEUNQ2zJzhddPZGyyu1YDeEE9xPJ4olIgNugjkbszoS8+b2+IiYyj4nsbRgg7cWrjt8QU6
LP59volQCLYneqRVk5nLM9WYiolmKquS/RPdw+d/Ou6+u67BSPwXkvWNUoIiqLEaCHv87NH7yhip
9xsdzsfMedc9COq6I38ufS9cugjoNi0Wy51fPDIP1jRAFzdJqitEQz9CYU/KYqkAUHsB0U1al/LN
7ZphVwv4KJcimU+kHqlsE+/H3v1eA+/vZtYPhjKX8arkaV1N1P4vvRvM/LKFCnncWZKqDNgsPt/X
kZ6J2vgcOb162N4GAh7aGdI20l9qz0wALXUhXzgUSpSxK8hHzbcH3igpaCGrqYMNoBW4xJjrGX8g
5e3us/dRWUFbiorG22h82bVA9PDrLdvhR7hZHoUpmZkoUnMMU8YlP3oRP0aS/P1g9tAOb+vjOCCl
gwsYre3qMktstGXNLIb74cYGkFoIDWJuIXphIpxB984JCNYcE75+NpKPRGoxkbVhsLbuiWFyd4WV
Yxbz9/5saadj7xoICvp2PluJh9YJY62lLsx7CaPYidmiKrpbaNrUvyaLsiJDYCHfZ+ptcLSPl/dA
heP4sW6teIs5e8u3v7Io2Nt5Hsbk7v2pMDHeUdBM9R+H3svZa+fFuc6vfNp/OHha6RsylH236Gj4
6q1pM2zPpXxoL3+ng2+3ROMCxXuRrdPJ4yVff3/X7CtPSaQMRuyvBBWaTIMFQqkv9GBVyEJ1ulOx
nAckecKGSzALBC+vSyW2mqp7tqaUEbklps5nRiJ28+HmY9rlL4D9tk+Ly78O+Jr+eL0dX5ynN5Vw
vzA2WiPZrzoHj2BOqodKEBRE7Mf3zhwJgVez9Xy+tZxXQa0vQW/GQJaWeEsjcDbuV6FiXURCyHZm
a6WZg/hi2DMXRrl6922WzA/SPnXH14VrsdTYl3pdlKPOYW21yY/AOFbFlWqQhgAilrjSjuM+0JPE
3h0Idkmf8u9i1vmc4ylwU1Ewd6U9DQIr4LGA4SxLfwxCHNBE6xudd4L6UwVPCzghQQHGO+uN/c6p
LCCS55gF8iYjDyEn/yvyWxrJhLR8fXsFyZSiY3j/w4H5LdGASjRyFd7cxE5oyx0Ib841bkhYPlvu
u0szNLH3OAoLIg3Gm0Vuk6S2GrtghBlU5/+idnfo3DFAvvr7zBzpT9OjJQpbezzfnScDWZNBQtTc
1HAqiRXMhoOlf4pOxQdrPDcpIlHQOY2b88TFGq42HBFAltMHOku68L+VaDBlfRbGpisJgUAJoP+Z
8b1Lxsvj1rzK82GlCEWZ6NuUOMpuee5I5gf1kpFbh3raa1cppAz7ffsiOSkeMwrfhSU0S5DQh773
gbAztmnTuc0Xcg3dZZfsWLwT6cxIVaSZUmXAlZEcBALer6uvhn6QXPpfXfiymBby59YkJvZ/0lTy
ZbF9hG3bi+6VmOvsIptgBqEH+uILWygBg5ghn++B25cETWbBNmhvYdGzZF7owAjCajhdSQJutB4a
VcKrwlUtpIrlGlj+LXKFjxXuLHqJZLpWPFpDCQaMYx1Ue18ghc1l6EyWZBc3FYMAijNPGUITJqxY
xye3fIrre5PGAWmIWEjMgwFGS6VOdzDR/llMTNHq+GIidfo3GbANtiSfvergVx0oGpLqRKMKiLj6
YoVvyST9cmqb3s9rpqS68sG2SbFirT0b7CJjsjFRd4z4I+htTrVGOVxEMnVt0umnTPE1a2ztRtQT
AZr8LVZT/gf+HFKKDhTyf6ynKEG7PFoBDBqouMeZf1+bviMBkMortyY1ZU/Ms7L/Ltgm/HQQ5RPj
s2Bv9mqOyo3eTnTxeb7i4IFtaXodmzLkX9oBvFjMS1uLqachE+Be2In9YwehzIEcS7uXtBGOaV7n
G+V2IHOmhoKHpM4DKijP0MgItggoKWS/q5seXIcql0Myg4c9UYYmNFCrNk5Z6PukNOPtLEj15do6
iK/seBDnfka1erL4JJn+nHsMBP+RbBOAXG2sENjHJUQU8U5ntwQKH9p5kck702YLyOsOo95RQObi
ELr9ybLZp25oW2J4XpOs6gfhenlONAqQs2w08UgQu9jFQV2a0JEmyfhxrFKMawJoE3Twtl8rx6ZW
dpfaA8mATBrtxeR/+xLg29jg0XwMIod0p2qrlB7zHsyoSn7ZPRrq0afaZ22Q7SKjJdDgsGet8FlL
HR1aS0gSqqedWBtytNB6pCWVEcnJ4f7RoqaheYTYhC6KfIqgO2osRuBJHCwkR7qoOzf2i62dN1dc
9SF802iDr0jXqGYWf61wHttVLocmLD0ciVFr3K3itfBtMd6xQDmgLW2ssNxTzsVBNbCoKdQTKC4a
fRbBlmGdTatVsnGVd/PFP5tDlzuLe7q87gIrKmd4rH/mydPskPz6z18zud9EBfiN+YphWhi2hMW9
oZK1YTB8Xz70J/p32DqN7OSGYXPXjXpeLHgUVQ+CN/QLo9GVrpLJoNqzKrkcbrBQvV7AcM2eSVqP
SfDPs+vdCCf/w51fuUXpBdYb9IM/NYZncsYX56VST49M/0RFar3JbF7Ip/a2kotq9/njoz2itiuF
LioXbUofp0txCY1g8r81SEKcQVipFgxnXRCvz2uEZirT5ggFrrQKFAuozc0vPEpE3hxC38g7RfyK
6o4kJSP5+w3pZyKoyM2rtQ8uFVlSV49VslfRufhtZGE59giE/l+lGESidypCYVXdThy9vjoQvT0i
ht042+8k5HRB8sEaT84Cz/ufTMAeQy22cSCuFuf+heAxox702zpcioMXEotbKYvI6WIGBEbkpqe5
o4sGCi/JNVRAYVJMDaB3kn3jVprTow6XCMX189ZL3H6Pq90NRnfISC9vddQgbAylTRJmo3gsQ0JU
7TJcXEr8GQAtTVmOkedCWkNufsqJkDFycJPz/dvSgBwR4+FeDrnWcP2iLCFvLWkU5bIUEIb3rQZp
rfuJCb5qLZY1yGYUYwPJQpsOj9UIwV5Ht4yd78SaycbSrymlQU1cJBdmHow79B9tRbukg+9Szj6+
ATzXNkyzeH6hx7zTPzyGg19sZrNaC09Hl/9qfjpeSbeWOdrXXA/RL87zvuWnFXxuorsojlGFafwg
DaBpIhwUfT++xFxYtHC2DYOtnjdTFrm652bN9nTXj34z0OGe97sPUBIMNez1J1xBu2TEHBbknKkV
tRRSnDuGoDH1Wzs2iwrAFJ+SH/XpFv3M/sG18e4ak8/dpiEVciFMoQgXaohStih6dL8W3WhQ2Llf
uoxB5GpmBshYL2QS1YF2cUwKZecTYt5TwwKTxXWDnb35NijIE1VwPfq8As/pnrK9p0v4qNFiiD74
4z9LKUrZxl0e2t7z8CVRIs9Mx9UbbZJQR2wGM2FMcrv8yhek5/QA1xA31nI5+8CBUdoQ0HBuA0KM
u3QxSFY+agw6QNt1unIuayPyjcpSMW9izmvVp1PATejQmlQpSJBILiRUx805r+gmKASWYttvJRnS
aSnh2zv0kBieQjH2XgvOQSxVSphC/bHKr8HXwSPgb69QXoycOvNfhmsfO+isuepmmvXfQSufCjQt
4wdjieEV42j2bUZfdrDg5lEivEveJnP+Zs0ru7UZLw+/qYiRNpEGQtkEngSNuVnSzx4xZEFqupQJ
UicYxuuLJHhC6vIJVm3ZDWSQJPVUuVHgK7I2c0bpHq1FOVqClYoNo5/qMWSNJPLAhdzjYn/YycGH
rkrU0OYTDaIo78ArdlvfEWSFDzdPYsQZStfhug3XG30jhn8S7f4sEN6zh47CG1/1AcFJmVxsefD4
Rp1jbKq5HeI8XzAjzB9qI9hDvbqIkNQe4t9gcANtGDC8X2DAJZm08qkdP/e2KtCpFEFc2gocZMUF
yz6MRNczXSLukYX7TjO53R77w3MNjhoDuuDzjpGgSn7lNPHIdEh7DCXq8Ba7Y904OFcbLKtvyYT3
BFuQRIOQ0J9aSOEeRdQNPcF33BGCHBwFGgn5RSM408hnbrWmboWrrLQr2wDA0osh8Qjf9b9uUTYR
7gwUxttb8/WyqCRjFSM4fytmQEAHB1GCSF48LOy8ZzyuVFYPy1/q3yv5971HqXhj9Oqhh29es5n3
BnZLhbQaTrZlzJVmkf15oETIfDq1yaQ7lACgMzNGIBqSAG+cy8E/8DSAvGBhkzZ/qkVcAG8NfhA4
KJ8uocBWW4FH4jA9714/19drRZCLVJGsdjnmLurBh1X/Ze/0sgBi+bS33d/S0ED5YKD5VanXTIOc
f4BEl6Aq1daX5QSAq6kSH6CEdRLJdWjfeT+JB0rs6LbMSmq2yL3NyALv+nUxXk6ynzbEhtAWPSjS
S+AX2krNYQ+lm/Wops5wTZol4ss8QwILaM8FG7UHNbqDEvdI8DVpQKU9QSX0cynTLjUKWhghLm+L
VFoD2WVaTys595LxpumaFp9sQHp8soKlP06HzhKUvW1ENOijxcd5lqc8F+PfHrwixr7fj0ML9v4v
DZrEXJx3gVlbIAYIdGZ+PtcIvNzTmhOZbGTNrIaRICfrIxTJN9RMlr/vjOFCLOLVYmWn1yidvTjM
6Epl339bbafhOB8FBNR0y0WT/UB9B6na0Lrse+LUxIAFxwzbDO6XWkDXB/XIBQKBCb6Jj7SfkUNX
C0r2cutLQLLx4+HD6rk07rDULK4qnUBDnzZ0yKLMJ0EN8UIeuGKA6Y4JxB0aTGTQVStsUbmqHyev
qocP9F8a07YRdjEkZaNFo62OUlVa9htqTASC7jM/+1pAyw3H47P2ZQd+Ie66ZDMblTc+7ENegdSz
yPMj1E83mWAbORzTIOzqakL7p1xczFBEz/NZyIUuOx2z6GiGZ5dTCTitJMBomK0bLY9Myn2LVgjW
Z1uMhREjr9Eq4zV5+MCm1KsGhZ2lCbqEGtb8IpCYegLQvAsQl4Fi9vaKFb/8vFMXt26CTxnX8CQZ
HzbAAuLhmGlr8hJvz/KA8IrSIcRiZAFIybrQIR/pEYHW+z6GC65VccWcVE8xxIp0mMMpJQ2dIJOR
DLTYOQTXVER8nnt2R5XalMqGsZE2xxQMTZL+M4mvkJpT9LbgetmLCj4E+R9b3ugnjZyqpFrJtC4v
egVwa+i4d9xQa1BATGiMVrIA285r0gNHCPTXQE2n/xBbOx2SpIaBhNR/+4OAe9SRswCuBUXnKVzZ
J63b8EB1EYkmsTeKCnkU1aznXx1tz3kjYV0fYd/NEoS/o/jIeARjIzdB7MF+8oxqVNV3cP8oFV+K
C2aBNShqv+bKpKjjms1NvugBB7n2lPzD8h/1mguMeKb1Fw3MpvPNkXyTAuiZGh4vtg5faW3k2wJm
afsDXveQv4DQRFWi0RGi2wqt93H2KXTjY+5QBfGlQHInCVk5RxdgjGyDDlrjTgW87wgYBEPtyjuw
hPNxvrtg0BOSQiye3T42QEWLod+/5xatZ4zvCnsfXzSFiNsg5B66UioAR0vgWXrzjkaKnDWQPRuv
XCBRpGue7gEXQCIed8HgvZp5U43JLtfPWYuCXRmbkjzrZxERNzdCNj8yyL/7gkFvPJcWC/IAZAF8
RRteCWJ9La2sCxuXFzKsesQa90V/4n3lzI8b7Ak/Z57/OOE2t8PpRpAmpu/ru0U95nq3UbM2geRb
hgHYiXn9XiC4dwKuZqk0P1qlRuHpIz2zZt47f2TyIEOp3FB2nXIujFvNZU8Ddbzgjyd/yJs2XBKf
fOlza2KJEAEvIA4RGtkA9/3JQrFiUOBIaPwNJryPyp0P3x+bZgRt2PGuTFAAtb8M7bb5/KW19B/W
3oeryHhftagf1dlLpPW+an/1U2BniDwFEfxtkgVt5xAS6yP+QyG1Fwb7jlG9dYuZzzm8Da4e5+B3
Z1NmxNySnmH3+Kq5jGC3qJZ9arWgGI4DWjJIGlrEE+8m8QSVKgBEP2hPcYU0RaNJHe7eRxs2Of05
w2/afZGWOkxuO0OZywlepAbNnYb6xPs8mtRDp4Q5Jyt6SRo7OsRyzLUgkTLOJQQsNvfAYMp6Do1Q
B25T/oiYemFWqEt6LmSHfR0/jmTc6Vl5SHcAfEbmoXU3cSNv6dtJd+I8kIvjlyq+ELJbTWOIJpUu
1sHtl6rzVwQzqwZxgBP2K/Nl2uQhMNJVAyRQr96qZO8AnYHCkLP/4b1PZH2JLKA6IiXkOiTbgTtU
DTB59KMHI/2Z2RP4VoSh+KPNl8w40A8HC0jOcogB7G6gXOh/uuzbVhxcajZvlcjHltIuaOGs6AhU
YcCJQiW87A83mmBvPn47r9QjLQbDWr0NKMFwCN7pZ4GmF2iJmS5C/8rxYH4/ybvAyff96T3sZNCG
mQisEYc9g1DJTcFusSRBYBYv4aK7vAPKsjfR5+KZxmUalp71xqdp8Ab1+SxGSR3DqMc+HdgMX5SW
K3bFI1hM+7H15ARNxzMQ2i9+r+qfmyalX5o9OiEvT0hLOUYCJYBV+M39w0ciqaame0UZkJ9G52qr
z64lYW/GrJe/zJ20yD8kWUIYMqUbO9p6ZmrHNOPY3f0VQCcI9h2gP3zOw1q9Hg6MG6LhxoPW/o5t
ouhKHpdeDrl+PjCnHHOhOOOdH/NzpXiaa3PwqhBoaqPK++QZgyomclkargFgFWmeNJ3O0CYiR17E
Z/6yAeKu2RIcMtt3nU0TEmO6uqcwRWpMFRvj9A19/OIQzcI8/O2DCOTuSQiF7/K3Iy1sbIkS0rVG
6tmjNjC0jtqM2/6XjuSmQ1tXv95HWI39w6LK7ee6X6SgrNFp/TNOdHow7ArbHI7c8fKZDPpYDi9U
YBmF5DoPZjEnS4lLGXbW5LBdel7DGuc/TPPuyxMpAlBc/n0YGssjYn/d0NAmxtv1/5P7BxQT9V2d
I0B7FWpXCOj6ja/KoZssOU0lXJ5b3MIKXLcPA76MZ+gniFPyP2G++XTXxbHwvyKdzax/nRUxqgOq
Bokt5ITrdaPfkKDnYKoeJZXa5KeRIRXeIVAc2Ht5Ygm1+mY1ErSyAgNeYtYnyJ3ESJ6x7lq8JNeG
ugJmMYcX+nLSDrTulFICzbTf1SgCpgxFydEScgfgQcN5wkp8srZ+T8rOL6etzrduK1eiHlJEgUyl
Y6aEWaG9di/IO71C25uHmnAciKuBmk27H/YBQP+lq4f7bx30S8WG38rmYN4DnFMtvNqAFlcXNlpI
hakys0X8/gBidTBdvFzB8aSEv3yMkN5p8s+c+jp0XxB4WdJSxrFpmaeoAahkBiLdzddHgTkRw02m
fhHUMvOB8br0519VKe00NKC5Rm2AFlR2gaRd/Kb/+vpUgUi13KB+iTcgTV5/DAdtWp/QTidVtavI
UaEln32q0fcC2l65ojGZ3YoZUkUyrukq/AEDQ8iRdglQCAJ2+dmiKbnr8bd9KR27wQ4nvB6+87IE
61RumoD38Dn4TEX230M3kA0KBFxteXJwAzWxh/Vez01T0JaDZttX1iEsCPLJGTVuJMMCowudQcgn
oz/sbpIkHrExZ9MgeX+DPD3AzIzU22S3hwpt4ZfEalUXj/z4BJut15EDhKV6ddSNn/L+l2LooMkC
HyV2apZ0oU3ePt2ckLo+BhvzpF84pb2qJIdjjq7Nl8atNfODF8Zh+xqauFzXAV6VVl9oDflTBIai
DpxTpyXwijK2jFUVoHJwBVcxzQQFQfz6JDpe+wUWiQaMLI14TyBCQ37aNBeqITOq7OJQwV7ZuFDn
8KAiz+pSJpjbl2DJZvua0MqrZ8oPXWg8wU0lfaDVsJsaxQGjhIgzy10RP/562Cht/DeUWq2c/p+p
cP/JLdTiP9RNMJ1pNBxv7fMHilsd9vrxdYPC9j+gHpF0OS3CerMZ/S2CbWd9/nJdnEeO0apxBXkr
Rb2/ZntUz4wjexZHxskVO57XI8xnnRvsWkJb76QGEqwv+P5VWddrdNKw2e01QoNRwCbwmMllVFdQ
0g3kT82FC2QiGqg1FZILKcRJr1m2nOA2K+TwJCCErny5qyGhtYcfs/JfwcOq2akGVkChP9kY/aR4
DpxIt+bjz5cpaF+7uRFq6qFnRBNYP2fiBOPCq7JZpdJQH6Nudg/rbqOB60d88wEnp28rqm+puBK3
fCNeHz2sIlRhlb3hVgK4tiHaDtmYnhL/31m3yX1ytrMZ8oltFfmVLnY4t84oQqNwYviTLJOeJu+u
ZpAGk2Bc6dUcG/eE+XypPpuQCuZPUzaBGCojAcFqb4C5NzhE3sAES9H4iakT3+V4YTXLGlQi26PP
IRCYTU75ErjKIpgjySuBvFTEEu8u6RdulY5Ldtv94axrKHwEMscKW1Uh0GHQNhG7YBF6hpDPZY67
+c1rJtZXHTBoi0sT7obzKJrABEtEee+iZRSFDp3iKu4D6PD2ZMbdo1cZJd83LiAWU4TAtP+ejFTb
MAVJ/Ghst1VhVsvuR1Jpnze7AbXUe7/SKDmEGCM6sWLuBsck22BUYF+scijkErFLaw7NeOJFNWVP
fgjQ2qxPrYrojSLsWahetgSoNJMaQgSqp+6lkYinb2xGjEGt5zYZDMTKF6SzuST8rOrQLMjZBnrP
CcO+5Rdf7B76PeqTHywj//Tm0UlMmvHQ1I3nTAhhn7fNZ9Eg8Qs2GFTHpXhCUlLGoRg4ILd1eBTW
UGXGxGYU2cCkpcOYWs5UxDLCiUkp9z3KKH4+61vyidW5tgIdV+B8P929NIH+CxN4pJFnc41SapPK
K5HgprRsVH5KCeKwl1Q2B/ktl8ebhos/BzBWwu9nu6SxbbuvNTvj/dsP4DHxrF2KPkMDUjyZVYcu
k513pZsIU6w/dl9i9Ekj40ILbpfXhMNFk0xiWm7iQyGlAOOlwwr996wgZ2dkm+ajXF0L2Uk6d23g
4qLNvZOYjgqreL5wRnl0Ru+OykBj2r1b1aTamI8Xuj/dEmwRP2KIZ8zAM42KsdzUTWQCSHdYR48S
auIo7/UpNGPMOzAPlMH6I7exLJlpBt15/jKzdCzwZj0Rb9PEUbBO8jpfVvNeZTlmlVcHZ/ntlGUz
s6z70ZLeM7vPADorli6ArDdDAYhoS1qlXD7W4l+4bU9j2ClNyhSIHhYimI5ecI3/vX1OXHznrdjv
NT4pSxtyx37HWVPKibDbpuTTKXzlUAif3GuibNRyk+V8UqZxmSkgvl2nyhgADR82aaW8UmrGv5dS
sYBEtfMlZxwuz7iqLkpCnvwmhplcT6yaT56FBJipS+J5H3eamRZGVDZdXZDbUcRaumjmTGbZ0wRQ
wgtW9KhrR14BlRqK0ytfY6bNfNX0msXfIQkieLh0BvmgYFcqQ9fjoxGR0FYUVtUNyBRn5zPBqyoP
spbRnPT6pym5Dm/tf2S1mDbzRGTK32F2lKYyGcBxEN5ywl4Q2gIOY8ggAFmxnvJBvqF5rVs/De5/
j0bhuWZ+UeX5zI9atSFJF/vbbj+rhbhCirsuX0R/7g7crWiKNi1jQkq/pbvq8DZpJm/9PtktC676
ZreSrDgX6j6EBXN+9vVw0M2EXXYaI8AGfb15A9G8/8JP/8kApXTNg2+g5QGV9Tu4bXPSXTDXyw6D
h1fQaIQ5D0ZeJFukIxK/eLyxk4tlCzpu5OgjywbG3r4H4+KAfpLfhH8SxVxNvi/eZ2JnAdr3zAI5
cw+f6rGaTWJHXdsWYKQrCozkUj2sbtq8q8dbgwI3ImBtwl6HZJeMkYK85LqQ2lIRMpD4Ro9BJHQx
MRiEBphywLu5O+5nNmb7lZ5HOWDasRKSdDt/HWFO8+ttyrfRf4tzOxWpXDxB8iz16B4VZI10DYMC
ETV/7IgIe4WNaXZwm9g1B/Lr8jen0IdQ+PyLpH3WAXIpPf8Pj3d1OKeHc1n4BCzhNIwCVPnii7GJ
cwV2TbQGak6Pt0e0x8I29NuhIGBzXITzr7MjYckkbGx/Ijmy8JVaprFb6Kfba8SnA3L55OSpkAJr
WLtjIPA/2q0J3ZJIBQaGAS4y8WPdBPR2jXRBdjc0eUBBSy/KiOWiVVEB771JajEYHfABIERzqLm/
f7bCTThrhYZpXkd7FdiKZPy5zt3+srbQXSjvBBZp9c3QlrvbZtQ37HV71r01L603TVhxjJyrR11Z
qKi19sL9j60cIxMCIyXBoZ3RJ7U42ycdOpEj1FTVF1qdj2vIEC9s2ca2Dn+zf4w7rfPcJrTfqA0L
TIz/fDqAG61Ky62GKsUcg04GXdn9Kc+wNeUuqp1e1rvu27IkddYt9yX2ih1cmK4VYCh/rr3T7E7D
NXwbTUTwCNcANCdm8T/hYgg0uLzR/ov/kDm1PSO9+GSX3ufIn3XVRZR48l1N1s3MLyF4I40DAGpn
YcbZOHJWTierlDKA4SW0Y7Qj1ju/tqVbv2FeLqb5bzbV7d+rTavGIahpFEfjxcQ2hKui1LQbSR3Z
2XYxfuORMr3Mbw/4DCsLxydAT2Hwyp+G7W55RiAkpiIecCPyGLWpZEE8aHxC9PR1s9ypI4HEWC1Y
gnoa71pOFfRrimF3xS1zMzJLMd9inNVOxXRLi8/rkxVVMe0SAIMiqXJZgXhv6cYJYqFr1qH0n4Ty
Jmv1+SJUmOgISouyhE9cwVnbVC0GXJJa1qofhUf3G94mdKawbrgvwZ+paloXsRBA8ZIdU+NRby23
KUYtxzVitrqSfFhxRdmi/H9FKBAZTeD93VL+tBEPyxYY3/wbl8LVdNc4vLDND5HvcVYfSUu4Seol
w59lz3/LV9qNBRlBJZLmIdMDG2QgmCosS2oWxb2OwHMN7yFwQUVEFQrP9klLHYDC0Yaq+UOAWb/y
2NNtvlVekIvbB6J7JhUMMIbQAvAdmBlE0azlCO0fG89K54pIs6NXTfMEyvPyQFlNIk31GrK/QutC
gFMiZfqfJpLrEMpsvJQQd3l08PzJcmnolUIs3uFIoLO0/u+xXtPbsZ0/BKVDqirWM1BCB5YB87Fz
vo9B4S5SnBfZfSGIoI/QhLOQNirYGErZjiuK6LdC5pJvzHxt/KNGzkNyf27YnHvWVJDucaRC0kIm
iqjAMgoSoZe3xil5CUNPjgYZUsBahaqUQm547vYZ6NnJywpFqrEl3RxEeMa9TnxjKo5iG8bSqFaK
K7IikOfTg2L1E4J6sDVnGGairiSntVSR5BQCh3HNbIG5imu6N8b+WgTyuEcW2UrsD6/Gi7+BK+MX
jaF3ileRj2aCdNGVkAPZDl2Kkf/xAKeivMvhBpz/NXmkLiGSlExU3jxZ3h0G5pMKVwcj7+k2y+hF
/Z7KoPENO26odIqRZwKYhFbMkSWJHm9swszcYMo5Proj7rTV1UWRtDkrECx+kl3XRB4G2MG2vgDN
asawEys8XeeLZnkYdl2h+ESue6f+vTpr+YQCbn8jxnu4je8wOsVagpY4IAoelHGIFLwFah/AqEAW
2Mwwt3H4Sanuh601q/KtzsZnjeYzRsGhue7M13DN6ARdK+l24DxODDrKY+phU812a3Zaz4p/IhOH
SU2BJOwLW9gaBrsJu1w3K5UC/QwmE6MUkaWk4DkYm7SaxlN9UYlcZ8Ne/3OxQ6FiJNe28JrrwEGZ
pvF8dvrDPSC4GmB5ZkoSh6P34zgHTmFvB0cCGD5DBJTJ1Qr2jTriXmNrd9+xHC8jUsNnl80dP/6U
PCKTEjmYcFn78XtwLWuYkVoec3ptOHy4AD9oIS9WActQ4kN95RVN2lNq+GF3BvHx15t7zJ+GTjpx
xgD67VKAX+98wx34S10VVFekM70PdgjJcKAJFDHmO9Vecu5tvZpI5nXE64ifpH7s9bdZa15j4w6m
5f4OyjG/8cLOcE9aOyeCc7fal7xTXCyN+6rwV0FFQlRmsFEhcIiPeRd+qglSibI4d5ypVx3CcFjD
TPol8h+iXTYQAASipDf014CJUWVVG8UGS1aICQ4NBf3rWyPUoFT9mxtOL2lFexQYvbC5sCO/mD1m
Hg8zAfgrG35YrcNTPDHvJhe2Tgeg+laLwUfRgub53/ucCXZnAF386d2twfWqnpxj+OhxQaKdp3wA
EQjS5tl3nIxk43AMhA4hJREFfph/FsoYpjH14Z3SKc8JEuIRGTZCnJgJyBrWbfhqiVPUvXPJ58UB
RAnl4iEDQedsS2Jj4PxrebwWfCSvIx8a3bxgGQLZLg2TbugbUZPUMTYgVQmOb6upD4OPIzmMP5Yn
4Am3qfg4eFESA/5kAoSiTM21O32VrHHAYpyJae0N4MIZpg6KEZTvoK99GNi0JFAv/qobRghi3tgV
rakVlmeso9G8fXYxCEokpW0j8TEKBVl0jnYGN5Ug17ryU+euNvMbgg51RtCqu+8uqgwZ+MIsdtqs
Kk1siWfOXyCD9v6G7DrwWYF+hOuslErdEWSSApLQL/66aroyHtlXOItW1sNvSSV2x2P146+ihifI
8O/nxTpx+KF+MPMrtU0Lwd3/coYBr6QGkgF9gJc3sYylPZjbdEDihdtWZHqSIkqbyoj2OrZyBMDU
vF9hbpEvW7lHp4iTwB28jLrwyyw2dQcqxVqo0iXmbTLGtAE1zAmNvw9m1tr/p24qt5tsIfw4P0S/
5qIRNcAvKVgw6v20jf9lNBKhwNIuTaS4NnPuAYF91shJFHlvkvZGrXf+DQG3OwxMM94RgmtSokFc
ykI8pAzD2V2YFY+vuYlnhQX2230Z2rMcx1Ecj/F5Bm5ACVLbfUWAkfGvlAisTRixgt+bASecT0+P
Q5o3/O/xgHw+JYMBKZ/TRNeJgZzRYz0j47H+fmGmT9SPJaQt4WOJxK76oATspEmrRfp5PKTNNZWC
4Mx1SqyM25zmpTy0Kqzi7ZzjesD6c599IiYbJZlgG7amXAJ3Dt3Xu/jOHXfOWmAWHCJmmyjxsdGs
l5D32DDgaJ7R7WGTrskoB4HISw0hGRt8kDcuEv8baDzI3eY6FT7CpwLE9fsnqsPzFWMpd/+1fkzb
yUIS872dXKpV6UEwyijm4xznNhKwVzQ1paFW9yFh5OdNfs0HeSzt0jA9P5rYuppGrfdQqRCMZjBT
TTebPE4e0QBtY4tzLPfYkekRIe8eGMTr9v9vbibUB6I9UdePTON5pw6IJh+yFn871EpF0NjZZeaE
JhYYKExq86MP9Wr5odnYD9g7ewPvlNvQwFcw+N2VOrUT/6oK9rNGfFahuH1k1/w4F2xUIdCzJvxW
evqWFcxBva+2MHf+wku228SSm6ECUVnQ7aWfP2UT+3dwNCIGALQlP8q5HwlfrQdgHsKtaAH0sYQm
9KlSneZoNqtzlE2GPNoOvnTuE+tagyy+dFyalES+Y4TTdKPgmvLUSNtOuGQ1hdev2ioYRc2vXgPr
hUJBWJj79V+rTq+X9RlwxsXENreNwbkMi5iFFkfHURbGVgUmHcY7mu0A9SK+WGHSJrxGAgxxe0p3
NiEy2eEf/JFxLDRBAlDOSuUb3n6tTXxlJCaXnI4f5b9F8O2paIibUB2WnwBTOKXhgfuSjYlsVBh3
nCPJUd7L0v8TQ/JL4tV4DqKHQcJxma5d//GODRLySSNVsK4finTU61v3ngNDRTbG29hgavWbakll
gb84AgUrxXQ0X4wojGrEkuQ/HnjcfhAXzccvX863NKGhKP7HAcDmSEPxI62UPfNTLMA8ZG47A4Yg
XRXg/VVddhdRAdRGKeZlWeiWDlbCs9oj072omd37pxns7ZZw2XNtaplHy/KGXc+A85xBa3sHtp/q
CKRbwa12bzVtWTTIPJAIK7Y35hHHisn9eNzLYx5vEHsSEmT5QTo068n3Qn8pE6pVREnSOvMKyMPw
CiWogKhyQr89iDeH8K+GlTVxYvf817Uk6SIV9JIqWwx/nkimvMCRdAd3vBeOZKECURgyvtflS4oG
1zlI1phpYLFKaff9mVqcdwV8jwcy8g2cVW27kbUMUp+BRso+zSHlUOzgWTihSRl7tT3z+yKGsJs4
IlN2dEkHFG1zePnQelWsZnINZXo7mcWy6YyBHrRBK49VMXPwdodTzIUPzh58WYD8m2NKHCVF84Py
fbwx5N0owfWz+gmAwMDn4JzC/QDuTIwffusMezdZBXuVsOI7r8+irvJ7Utg9VUuSLAAL7NxkuwcN
iGIRyBKHSEDTNlULY+mO6N/Slx0vE3hOvgtMLU8EpV92Vg1vXGp8eLgQJxYiiog3fKLLD1iLUKH0
6qvlxLuX5f++R66do3iTYF0XO/Vh2jd7aFAd9q3eOWXN/LFxOgtb8RXBzAjtoIBq/5ql/8gWE34w
4hKNqJVG+WDbd63nr7xy35LJ0dPJMZqD/1Q5NXvGv3BDFRTfmvRBwQ8k08fKTA7QEbiVx8IjwCz9
oLpng6mAY6S/3IJXlgh+/g1kiSLjEcFKZm/VP+Rzsjoc64uzhFYDrOcNsE3gB6L7Npozj6kZNjm3
93QJoXNl5NN1RokyzIeFpeFVHO9v64gEQBc18ICoqDNNNzt5fwMoqyaR6QY8iN5ogF9abaLbHHLK
shovRVnzMLbqU72MmFjNvKR7obTO+ojR1yJqdyrrc6w8HQ7lOcxudhvwj5Kgi2VdGyc+I+go9/SQ
79eurun9mBQXNIoKTBoGQ/PMqSbdPp8p/0W4hQEbSR9GX2rDa4jsM5lnil0PnA04I2iOxgJvVUe5
eSmIF44o2hbw/33R4UfCgqyqe8dIGl9939LxVo8tcPfdvqEhnqadt+0EGlCwvC1p/FTy4C0697/V
U+pHFBw4pUNsWtOHVFMXP+/oH56m6r2puY7EVCTF3FioI+xb8Xji3pNqBCym6EiXXo98YvzpOimc
VdS6G0eQlfWWzU9BcniIF7dRwHtd/tU21WNCgsGrsxKFpvPeT6+VMmWvFKb4GXSwL/1STtD52YZn
6Pk//1JHBATNdZ+n6rCTxhnEvI5YVxQCqw7g13PEOGEM30ibZbssjcMQmPVPGNvBKXUIXTqI3N6O
K8eVAcqeJ8vPNWd17gWfwsNJb5Ug6L23OOKQB6e/LlVSDrFVta8J/sFg/YlaRXV1YaDrRG/HnHss
tAe4D7KzfsklkLhJcwnZpLaFtAETh4IE5RhDVWoVXq2a13aTFXqYExs8wON7fcCj+t9VxHzPLkhc
0Vr3t59sJCm/OlT37N2Ybz7My1fzUEYoGayJcFcE4JqQ0y7fKepErECTvUGaBXDnymY4rlJEehHM
IMRqRlhJ9IrE4DeFI9vMP1VwBfVNKIUhyCP18MOgJb016JCzHZ2rtX57ML5ucxMwrrf1964R5n0F
xsbuSMeuDr2u3d+h2u6hWAI8ZAGs2xBeZEYcwk7BbbKN1Q/ZkN0DV42xcoPngPkAvxCf77eKa9DS
pQRO3hbibeC2+mF3/SdW3p1Oys+RBk37qRMoUnDS7KTHwYBS5dEPk1JYoAPZ5wBm5AIZviU4ga28
G7cq443m71Kw7r+FzJ6D0J63E3DKQD5jNobJhmo+8BmNrb1rDGZlVDRTwTZsRBKFGCS7kmzxQUNi
7KQqrAR0cRc9q29HPX5BOlw2N2cxhQLSqpICpFtJJx0gNJIxKl2RlozGY08cwedtTSV9ZhGo/WX1
rZbwI998G4Gf+yJKbHO0BDhXHqsa5viyFI43DTazSrm9t3jlw0YHP+7qINVTfTudQ2eQBM1ql0ak
4YuiQxZLe/YH45uEQY/1tJF6c37tkYqbjqm9EdVFoXLtCBFwPFEOwJH9uOpEXfvhvpOV2NMBlG1t
vKsVd4YsfB3AdWSjm6MeAK+ZtFo9jm84sPfRjsTR7ukR0iE5QwzIS8YawdGzctMsVCm5Va1bA90L
Nfx9vTQDFH0cOaqqdSlwlB1/QLq+4QDIDMZFpe5pej0p7M0ESoaYSVBVTyAdNdQ2/S8db1g/sw3n
z2dceMyembW+U2exSpuVU9wUR4xqp2mEp4+DGvR0bqNfoANHL7vvjPqhxMO2xDvxRqdkXIbPs0fp
uFHcN69rWhAuOkOGB/WPuI0IsDcuXlsBkVqGHPcjCb6F9w0tAEePHiPXRF6p4SUeUzHuU/7ly1TM
h6YDJ0p48FmynaTBCyWgNDhJpWEN0w+5/SaJmXbVbJZ2ushnAxfhE5fB3wqVetCrNNj+NLJZhC8I
g9JPNKS6XtnGTGaPUlsGEWa7YhY+EWkS+dypNe+oXBaQ9xpH5GK6HRkYsLo6olMv1xuc5ucSqo/9
A8LrHQQVpL3RR3vyJZ1tE83yRd5a1C8o55pQ2/f/1Vi93eCyxb6+tKK3AtLpNPgvLkn5r8DAUeaD
cP4fbcL2VCgo00vv3elbyExZHK8ByWgH28v2OdGUjLYvWVSE7yxAN0b5ubNp5ZJZgUVFEdza+8Hj
uxgR5iBNANRuJt0pmtfCRne002Lm4kj1mRNeK13kSGyxYOjALM/9WrA0lOlM0+1h7Hu6sjm47jYl
HkFV5yr98a4GoT7mJ6rYD1YxgATRRyKIYa/VtFeUnoJinYDPEsXbRi2GtA8rUUhOcJQJYpzw0HZT
d4q+6MBA2m+CRNSzhUI+blOJphv/M5R5SIAuk2rUyKjiHcf9mhKkWN78BqbjP+1Vh8yS/tvuS1wb
76Q201M/IRodm36gA8/1jgFh82klP9zPiSrHUSPYWACFqcY9Co1O7TFtts3F9rZRIrE0WDtcfDaQ
eZHAbfdAqaKR18uPCDw7wzifStA3hOwE9B8e+lJZeqbYJ5VIo9guZeHHgkH9vH7nBNZePloaTmah
mpdv/RqOK99i9bRGzfCpc+dBT4HaSiRMoMwrv0szfGXVrxSh7+HCOvPh47gfsJdfhcP6x/0cHvFy
53FrNddBV1StSOEPjMlxYVK0oXqxUuwVN1Mgm7TjHkUDDC9UUOUdJ95NXPRBuB9Mizp1LC2VSWP5
EjhqjJEhYL86L7Oj2l0xOx9DD1EiJ9a+imhrm0RaGN8adssAfUmpa0VNfldz+0Ly1J2b7DbuFRMd
8jdyvEYJ9qFWbNXzJh6/3l4r+bfi49+myuJMA7wcSnSqP/qnQasDKuc9LGq4XwaloHOn1bl2vBTZ
BHFMswxyEQQ2nrAYvxuaLE2z+DX99pmEO8KXq4v8MoZLpDgWRW/aW7gXaPyF2taYp6rffRHpAR5n
O7FMvw1Qp+xrD8enLsl/TN3ahkKeWldF7qvlfEv7inAQGe7o61hDYFo8tNzxpSl5bF8dKaGHAQv6
ycKim1WU9SLKPZOcq4v2GoPmWd5fgGzHrek4coNGKE4wrnJZjJrroIy9+lZ/3otswMSChmDEFfPM
giEDkFrF5XetiMaTdUKBEIeY//+AZgiGsDK6TZawo34zdX+eOzjxKbDw7SUByXSHdJhvgw0PJ4po
CSaEYfxn0LRAuHxodGHH/gnDpfLIAAjl+ag0C0nAQpOiDtcrWbbv+S8KXUSyLzKUJAQSezMarcxn
wFv2Oplfck/daYt7S/+E2NHUo0zkJjCaRKow3ec0Ik0SAPGEs+SSdM57BKpP/wb3kwAUHzCIXcE1
w6gcW3QpjxM8DVNsQ1utKrmvNBwsIYZFBo72CRplqz1xqzJdUleXj4mW/zzYvGK8UyWDJdUvYHq8
DPsEPYy6I8VLl+ifIyuCL6yTOQwgC8cMgYEnUhdMyCFwDEyIVufb1yc+Gvi6uAW1BEdOzxRErrdR
RoqE4r8DKsupgENNuJTqOfd9hLosVuBMZiMYDSoZ+iwDB+N5gWSpvpejsqPb8utT4Igdgxips4W7
rJgiyqbbk4qER3T5ISSIibsH30mxkbX9D8JnEOoRyg/aILWeQwMJYcloKfnKdGxlIhY8W9RWZNZU
uxHWeb7EaSF47H0M8uav6oocNsoy/tN/wx0StHoZyTR5I0oWP29LZoQAPsTA6qvDGCMirnObOvDJ
fD2Xk+eIAaTOvWrKGRiOW4e27KM0UGk0vE2wvlLu6QOua4JsbVDq///Tc+WaTpzvmBvkeqvF+res
g+VXj8qeg6PDF6FWwv08EDAWt1bTqk9qpk5vvCGLY1/0zc/I05sXgd+FxiiCmjJJ8w5YzX06qXfC
hteO8XHAKHI6Er3AqdOM0A2dA5/CZKXpim8QUfTSbyj/qixhZ13lXNsTC119A1YXTw5cwTCTR5RU
rVpHhx6y3mhzjHceht1Fry/prYPtMQdyV0GQGcWJSYg87thqpmpp8Pc5M+bKCUO19KP8kKRjHkd3
16GTRoJLRD3gCFyox/gXWj1JjRxTe6xSMcXCBlQUZFudqPUGT/vqNL8jPgfcdx4l62yXmjeTyk13
2Byrd6R2qC13kaCpnaBG45WjG/5mRS/waT4mHMTnuJY1s83u/t8qB5EF/cmmiN4SGd8+/yYwuJD+
lTnC8W65YZR26TzvXZhBrbn7Mphjq31g3g4API8fB0VS7Ffq4Ee4yNEG78YPS3n52Wr/4XWGtAW+
domhp1JKvjVwxFkj5zKwyse+oWqvkUVEp1RCJcsTo1STrdbe939NnAK3S5IKVe9WLP+SbTeFbOn+
VLM0MBIamJC0kUZpaJ3ZyMa+avzEMYZbEd5/P7R054P6X9t/ohBwnN203pHDdio3WItCFp/a8dip
je56kKq1Qh+4zBMCoYOhKm8E8Q0EYSsYXUeaf0kjfB2hJGEL6u4a/Ph187iNy0wdxeOQPgN6jkMr
2Y8AUGe1W5b0EY9hwESqNphyM9HWoPHWDDixtYr3jprlbTT26kxTuwWkc0j9xCORl+i+wwJM6FQP
S/VZfX5wlqBr1x2kQ7A0wiyqAqlqbBfaDpdLTMNfafl0IwQklxwM/TGFdC+vOGFsP2BiDCwOInrh
pzyWaz2hMqQ8Ke144L+2IHxAmTKq2+8aZs+yMCNmMOVG5Sun4LeLV55aVRJPFUS3BS3CsOcd8Ky3
yrC5qtKdK4Zgz0aQboCV0x4BchDez3qnts3eOK4Fn4amgE1aDT3QhDugZNfj9m9Vsfw+o72RU/sN
JXG+/jPNIEErH/0PudKhFxkDi3WCOODDIjo8k9nwZGK69fIB9cSncYkxfEhhWA1DzXP8pBCduDW0
OLtbe7imKhE7pB+h+yEds74/a5C7BSkgYebxJOGoJWwfI6AjO2ms+w/NadzZRQ/LRPV6Qx8z0Jqn
R9weVdArtUZof9/OPDtu9LzdicYcUfZXXY+LO7QiD4aDhK6LS5lIDYkH/YFz9CoX28iFb9JIEADo
LW53VypvHWDRAbbFd+tfMdYu43vdTatxPP2UU+CidTb+c50BGQPldwymHGKaDdVFJsqdu5hGIVVT
/6PVMpdN3VMuszpl1lc1kGVlexKS7cY9pd8DDAeyb/L3eHrsM7bpScQpWTazMyfSWgXF3+4cu1PC
Z7kvhUtO3gjiKao/oVgsa+QDUiZXonjm1bgi1qMKrHZUMvWkA6EjVB2Bmc2U2vL9xvCqRrJ7rAAL
HVl5vjAfnCN5qF4J75gy70NqAGLBpNnclUkqzxrMORA3+RUXCcCABvv87IFnRufDS3BeLw7cpnnt
WlXyoAwDJn55+zTORn0xLHDFXuSCfnSsE1tK5WFFaIQWe5+KeD5MCOkJjIny0nUZHsOIucQvTjQQ
bewPPr9Sz69Z/5e+4isaJxdTKv1XuMtEmKfBUiXlKPLqJRaeDWmMXtPHBHITpHXKg91zOnhwEZn4
kCCZs1xqZjmWvfjuYe5Erhj0ahH/uuqzi/GEQqlC85zkuyBSlUfw7YtcWo7JsHk0BnMjHRvNu4lm
C2KU2aZ5w0AKRa86n0YykoPf6Hg803pHElKjE4XeJbdDSK7Bw7S8zIsvmpjlkr74iUMOmawgRoGO
+R8EebYZvECCbyxMymPahpSZEytGwJ0JpInKml56d+PGETor1YF6PE+zwP/xjIxmPIkBJEdo/an1
7jfglhEmvNLdM5olhJxYDyEPSf2P2YGtfuEhjRtiJXMAGBIIyXFZ2wfyxe6U3Tq7thUE3+VJUCyR
7RwVOml7Yh/FvIS2ctWhIHkZbDgZ5EwnYReYfR6YxB+9U7R5pNb5DZIsGfv91XVgDLent6VVByYo
4vnOUhNV2g+TvakGTIQDisnluJpe80r7HrvMuqR2F3KB+/P6traevdiOALOTPBzcIWf3pG4nKtGP
z9AGY0L4ElJjTfqvhE8x0LSjrG9pcjrG//fIqAJvvZnWkUwsMLWp9XB9Ux7y6+92wPx/EBid0Z+T
tPuusekJQYwmLGtnG9KcZMd3GXEgsGwHNsI8xaIayO4ent+w88FT3yhYHWUBmPWVHunXibLvnFIW
RWPVe9uPZWUOknYEZck3LBdeq7hW0CUlBZCZ1WA682OReP54Y4VaPlkGRfZ5a25pDQOwBmkKV2VW
3//V4MJtHzHSGbvFPtqHq8/+eG8HjS/j+IN3L5H9q8rsYOVmQCL//WzszCnfMnTCH349DA+l1H8/
H1jV12Y2iZTChaFtnoGJ1A64sI14BfRbF8h1yhO9qlF2xAfOTDgfS0DZMi6juH3vfYIkH3g0yMyS
DpqVgodSSmmnHNhE3uczUweKX03I5jG7DCsw6bCleXU8iT96MMlzwCtgpzuTv6+mgKTZRym4ZsKS
2WUCDRwz2OYQ4phzEY4x5vfTpu2DqpmMmKuS2Fq6D7BopvkI9bjpPQD8d+TxMWtweAEBuNU35EKO
NVRtalUu6SNsE1XxR6dtUoxwtf4IRZgSfo2He+xHwvkbUTgGYYTjPNxcZ4BZ4ov5U4s1s6D2/ZWX
c/LzVOJCMjEpFApMbEtMydFsM4qlWMKcTNFc82tWQT2ydWFejVRyWaJOtJ4mJ59J7ugdQOZl36ot
PR3FUhVA0aEW+Jh0UtBfR1aow3Tfq/cV8cKX8kG2sxha8gKvttzvXrSYscS5zldxXAZgPyKsH1QN
R7rLs3pRYSLK+4izLosGvgcRKRBDR2Evm/Z0r4ASWjvjqamoQADpfTkzLQNAwF1bn9a5tYMANy2/
3vPPN6w5/dMRna+4uri+PQx7sOrvSRgzqT+jjZYrB/x/R7YnzMnPsPbiezCNs31SolN1rCM1yXPK
vXfcegGaSZkk5VJCudHj2PzML0RYEMgH/cafkPfgl2UERg4S6m5twZv+s6H7jit14HokyCQKKLJW
gpa8EqXPswvDT2YNuBzLj+XhWr0zsNHYXtfeiZUD7fgFuvodozXpmJQU6T3CZwv54xyxx+worbiJ
4lfsvxBcMBCeJHNnws8ZKaJp/+bEjZN9Q1rqMpKHuxakBMxUEDrQSbK2Hk0nXHPffzqpZgErvVX5
0uK32cGHvOxQTdQZp34aacDWvCmzrXEY/ACDovQa+b/QneeYXFmLmhIAPVfdeO3zifD+8KycP72h
EdcmefkIk3mthF0SzRql5xcr5iQYg5jR1UodTcHgdCC3WLi0B2j2AmlRsQhh6nbvAnqivdmReUdK
7FwLtnCYkMB/hDBxHzAuUjG3OvoeoFMdsUgeP04FUwM19ciIG6lgC2b9pOJys9iJFgQ68OQx6ATr
xCXU3mcU2Y0Ap61ovOZXNujfk3zhzRJkVMG5BxHe1C9MmC1Vo8XjHhgCDUWJFGgSaKUtC4GXXvas
WBTgh2zuVQxPe7YzmKci5LhT8Zxn69XxNiaa2OrDuIqxDqLXnC/39DPsUQ96HnEh3uy9/e/VrE5n
cTMEj4oYX5PW9J4tp6rJ1V8YYug+QQt7h0rpzLVHYjDOa5xFQaxWSWrg2uFd8sK9QjlUilxLvhql
ENBl0fO+by4kIdRilDL0IVUOCrBpupOy4c4rcxBf5boG8GA9GxNNUK44WTsz58G5XpLNQUduR5P5
r9PRi35gRPzbPTRJtW5KOCpDpSLGGm0w5RXgx+zXYRcfJ0kf9LV+ixTExeb/o0zVv9FeaehxuTzi
aRI9qGhVHYNGgT+P+2e7j7iqHWciJHsUkR9iDN3D+Fwqe/x0vyhgtrUrdrAuomyju0PY0nMjS9D7
qByYUAqU2l5RH6bsVgMgD65saGuFCBwA6yO2PqnWGFOWO75PYSv04p02FK7Dp866pMfQzhirGLPN
WmcpILoTQzAjVYhbdjQC+84bydKA3NiD9Z0V2JcHeNqQZZcSHgwptX6tpqPpwuQ/KCgI+WHhdYbt
d8rgRcqgVfT51Ral24RlWyT5PNRT0AxOdSaRaLfhgCBim0ocEiHQmtvhmBxtt/gD9p7xT0spbTi0
yh235EBteyFt1XflrZWaPNzPpqxVytL1TxVo8cMIfz9GwzK1mzGk3bxamAz6c23vlThkic9V1I5A
YDsQQTtaI0wYluEbZo6S+f1S9IgPOrzvAehyfTvJk24hKQNxJRFYUTT56sTpcwpYk+MKQ1ZaMV18
SO+S885UEW7L7l9/euyNxzve5DnxbwhF6kPpQXoGxNLc4KzP6cCC3wTMsKB0KL0jHyadc21l1TfY
wQAvqMAyfPhwnW+bRvfgcm/eHJbdMh0DqerUjFRJwZGIFp24u3ZCiskASIxNmdSn/Xy4NF5h3Gj9
cDM7RNAu729Of8xsjCGj390CT6xiH8a4D04tpMpxQlaLKdRBjgxFfcBfGI0shDGQlfrk5MIQj8VC
RRV287+jKjDZI1zKOMK167fCPbU0fcZJGpxNlL3lu3+30OTM1ZDtVFcoLiDuq9Niky+56E1GuV3j
cFXlEFfA/0NOS5yF3eFs3M68f7mtlpOVXboOq4FofA+v9xoeZkfqsaVRU+ELK+5ToEKBc7xOMHr3
Q85QbDtzmcsQ9e/cDYBVQuNn+ZT/dtlNHI+SsKDdyMAoyQ2jzXoY6gf725fLCJaVIL8fuqcjVz/F
ulxH/V1RMndkDw8JjT7UUOhcQQ4J6pWP0q69921aCiSRXnqXeH5dGMB/TTLAozzOaEP9f2EfLnYS
iL3SLpanrzTyRRzlqYQ5ZUoRhfesh7rXasB7gY6ccJSb1Hgvwzi7LoI/UxqTBI54M6any4d43wJb
Ta5xXR5O4WIcNmvekD0CoEka0qUhgd+2yFKQrMj5n0/gD3zvqufhoDmBMIrHR7YBsHyCJ4bzvpXq
azUo3ld3nnNsCtSd112gNG1gm2jkfnJl/w9HN6W/kbyQ/AXsZptnupVBDVRi3UdPyUIaWuaAOlyn
BIDxOfgsj3An2sXLbTCOLRMGQBObMBrrfUFoOF9nwfo/IlkhMy4bbFBk/8qdAjqCsr9/eAKalEzv
7U290lJGmXwV53HqJyh8+iU3ZA+JgcDyBw/IjmvipewmjorLwZUokC1RP0yEzYS+aKBpWo4/ulJn
ktqp+U91anWxBfQR3elcsjXdRfV67XssLh8NPSC/ATrGIVYtlaNFZIrwM9n31EFM2np3bxviq42R
o22B4YZllyLswC6YUNGKqSe+a9bJawuHRR2AaTC7lgROBUpAGtxYspNTR1Rf67m9tviCYHiPhMwS
lwfg1xYbo+SEUyAS3HsJ1EsnYF+2GaYmaPkwsQ/lngM+Ith7zGIJxXJdeFvsQhSEi5nTejhtJ2+V
XIwak6Xw5k+85gj3hSaTa3e5nP/vhnrkZ2g2btqtiSDa2i7fltQ+KjimXrfmgZkUAnA+u/3LO8UC
3SmDgORb6bgUT6ggV26mYeRBqFW2L55ZNH7Rb8WkFbgurNcZ3MNQDQjq5/wj5MlX5+hkznk8poss
oHEJp878FyL4qCm9FYD6dy13CM0H4Z75u70q/zKd4mCQaO0A0cc75/3w9YOGzciGFiqs7LR65EGo
xqQRcJ5QpOmBkGsZvROJD7YWYdDBEjhWTqZS7N4gnyWWjvdxwXlvq6LAtPFV+XV0xK+Ilrfk5/YH
EOOZGwZO3mpgpLl+f9Nuu7TaxdAhYDXs1FSIQfBWjD0FMiM0vhjswitAMC0GDdWbgFFV43De5F9s
zI+8sydvH9SPttdIeXM12FmdOUZrVQqBswzrYxjoYsCsz+/XJ3s2bE6NwtfjRYsnPqcZbOnUAyTt
x6zlq5g7UMplV/VXqItaiY0aBe7dgQErhM3Gce9O4EJ/Mv9tkkjv6ZhCVCudYvYOAUkKdIpYWQxg
g9QtfhmZTllqtsPYqCJdnq9KyXDdMqU2hrpuJUwj+DsuhHDtunfFy868B39kKiXhSysoCHrzRAyS
xyMHe8UIuxmd5PGXWyEcF+7bXghzYPR1h8hKavuQNe6PRHMHBLwIiCKzVva4jvY/ZrqZWq6sEGNb
E4CuUEfTtGAtcjZ5NmuCd+fjTSjpJMk7703qi6Bd0wzxdMlQG++9L7OkzbuABJZjknYYk50ObVYT
vFqHmc18VqKqGCTV+jZiJQvFLhkCvO3ng9o3USWcS/WYSyvRUL2uwOO1YWNIE4H6kZa50C6lHmex
RGVs4XUxIuYIL/H4CxGRIGA8+Ej7+BTWq5v5x0Dbc/JQAennBoTm1zkOteec8oqavWHlve4VB/Nb
fyPYvTKUVWEIdNaWSp+ilr3r1Qd7HHymK9hjhfdEh2HFNrZyCiVdB8O/O/3FWXeXP58NyBUgZWVR
97kKqiVhHzwC+AoR9Mz+PJLHcNrwihQfLo4MdPvXT1bltXq8lS5j4ogzkSdBMlggcPvL+Gd1eILJ
p3KE+i/URztXSvVAbPtIbDjXuYi6Fg/WPYq3l9X/l7VSfDQ/3VF6/7f8wA9NW4NGdqDxFwatyTtt
YSuz8MHx0KAri3/lBPvHMEVBHOsH1FEz8cPEa8U//yTLTWaHNXyZJ2ezHRYXE7vumzVaEMywIPkO
koh1SFj1v0Cj3dR9VEsjPBqld9vrbrn4b7oDFio8tpulqlmUhVraSNV2aSEWKJP+q1CzWAba6431
MSpZqPm4Kp8kDr3FlMI0CaON7FWLlRElZs2wnBsErbNZckpHquXgsSydT1a0eTUS2HkAkdLit8qa
VUXzmhCXkkUUWYgJXfD7RS55MLLlKh3bbqDHs4hllzgQnCjicbq7vi7d8+bREEGw+nUiGRlTMqBF
xgZW7+X4/YPZ/N9tMWSLhbzFG3o8kOd58UevkJlksLpYtdQsGjQdr2HtQ7NwUez+q5l5BM02wvPu
YBMXvEVz175/xvCD7TQb1UlEUgLUXtu5v22Aa4PS+C9xZltHye0VEKpFFCl+RatSP+QPfXtpq4gd
kgzOXikeznfNfswoaKUnev/fhWq3Mrlbj0GLXfbrXKVEjrUyEJF6CxxoA8h6T/zrvd6UuHM2VLfW
l49Z8FYDTpFasxOqJizRVtmtBQaQw/Lvd89Dj+9CXHpDmdFVmst4nO/LAGfprOCWxGenA5Biw27h
0mxiUxS2fse95YCa/OArRGYPgOxbXXoWUNXOjRDuIYDU4frfI2Ysjkb3YXamnbFdfibnzzGiSXee
8IZWJAWx+Z8gELkic8z9twTUPlRsYHKkCS0goNPxRt9j5HbF2dDyvtII+eJa3tWdtbyaSwnvZO9N
Nc3X4BmievPXJcSaHdWC0qkVTPlO2oBNsRwG29YEE5OfyWtiBhrgxWprPh3mpUQkG3V7QWSjbxTn
rWBZh1CdzUXAcBrRtSw5KH9ahlSumrPq1U/Z7HFJprsALKm+BsoCqG6tDFCgzUGaX2bs7zqW+raT
utvIEdZH9LiUWpWIYU8XyLf5U5sb1F2RBDmySiX6h5kh0tcELVJYcTCZjuAUH/OMgC9sWs+RsuiP
BBVDhVIMNQhMXH7XYaERIQgN4kVSELaghJgur0CqKUUHF3zgiKF2LdxQIuqWAPw6R3ghV1h5WnN/
xAR6RLUu5XmkzOMQH1dWhs7mO064P35YFCemH4fGWmAnbER4m8HzJlS5PnL2phV/T05Nmj6TvNDA
5lJvVRcfb5okkyDRTMne5UsF0BXUUBl7PZ9Lz5BbQt4bw/O0PE2wU/UXBaQckxcvShntHN6UXMux
7u2rWP6J9kORnUdQCTmZSowXRKKVAYsWgNJ7YOmsDeA+SoPIt49E6UkzsiUsY3slq28Uvffv2fkx
lMW/yJ6TkzS6TSHDxn6uK9dNWEFlqU6NEfwqZtRKfTxTLHO+D6fNPqJxTk5oF2s9EqdHN5wWfJvn
PxRRekkSSMPlUihm9q+WsTTiWlryH5riBnfzatNcxn5w1gnczpQebANcDqERQfeptPLRtcvhhOgJ
AZ3FGRKyJLcJ0kxDYwI30fUU8GEb/evHJRrZD1SSR2fV5CvP5uKY35ttkIJIqmGWQhBAnkDmP4jw
ZS88ebG93eL5MY5JnO8xXTiEYLt6qJlFe6AHEj+VqXJ5NDFV0bWoPldv0vAg9sgAO6ZvrQFw1Wu+
h1omT/uDlvAIzv2q4vTGoCzw+BZjS5Fb22Ptswq4IzdJjSpodMz5saDH1t9/KGWPxABA5Gw75qg9
P/neHLgtrgKgGwxnhLzPB45Rbtr+RloijgKHsqMROXUQ4aW0iRKO6fyu4EFa1pBqXDVlruom2T45
pASqOCt3A6+5PPu+rnb6gbGExPg0waajJt+HuWMp96cT9ivIKbg21k6cadu2cDzSUjLOnDFAfkTe
5JPwMlCSiRCqxWdjLF3ueWX5k4AsCXTkI9ZX3Lxb6l4Y1Xi+sFGcCsP+JUZXEkRX/QbJquRWLcXr
8Y7XuhMI6jM27ScfpkdIOwYJWp+4IJWjIhBznck/6kum/Wfl+XwkOw9UtFCvpZtw5IaZ53UlgMgC
ScpRF5umMDfUL1L/VTfKa1KR2/+V4NEhyGXvKYbJZCAolqfYE5K+tlmlTWGaX60CFiSrTHju+ETU
ymDQVZbf74ZJz+UdVcpg3HyH/FNE6k92RSIuT4gQWm+lln0xmlf6hBIGSPt74FfGx7b0nlhMQbgZ
4FL1utzbijWq2TvmhRqsnzKg5VLul3p3smhs5ajRVkScjMohkRYIr0p7fmkg8icvJDHxPWRXEpN7
LjugLicehN3ZUMKVJiul40nsFgwe5S91iW88KY1yHbA83asHiRBRv9qPlEQdFm+VGutymEMcdTOZ
gee2dZDpZTArLJU2LR7Zopi+cPPgQWVSsUE6FbNypTZil8uCEapS1fvyDfKHeVlSlKvYCwTff68A
a6LAlUxQjpQ4qIHxcpjeBaQfeO3oKl6OLc1RnXupEehm2t5K5yXkINipSCwTsksIS+kiuOFzIdue
How6Mln8oXieUa4wF11ze81DclNiJvtBPtMT7pMe5sqVvdvD1iC4EPXZhkVHdIeCw7n0dHmm2XkE
hZQZCyo75vT553Qo2rBFB2ooEIug7XThJANMi55PAM02VbxYvFHg02y+teqzKKYzHFel1LuzuraY
dcSU8c+EF2WK3WdGHQq+trfmqZharaQiPR1zspOJESxbijWAXB/Dzfy4vi/sOu82u4wcbtrVhm+g
kyyHxh5kOjf17oM/56ilTfuyg4+AWvjiN/KhoYsS7TAegrvz7N1k1x2f2ad5Uf77Zr04KcDzDaIt
dWShXZb5LY4ASgrY8aWm6lZuP009coRG5yDoa++PdGHEc5GjBrKSdloo/tIMGIl1VEonETXKnZyE
4FR2/eeiITHY6mpomd+xpL8uVsEajyn/SxQCHKBOkyih4FDTsGlyg5GD7vosdCe+fz1lCsupQ5XM
/zYVJuRxdA9/VA4dFmkU/22UuuD+qRZm57yp8hYFraTuCwX5RXdxITLb3WJUBitwyddNfkDbxgle
k//ZR6MZ4qrKc/f0NFaYSUXtQ4ZvmJ/a84tap1gB5xerJTdStWiWIKHJ7/YIPyqTDktTMLzc/pKn
LoTok4vUE1CJHO54eSaIvX2gtnqArW0XM9ohxJEwHjtFM5PBpDynrUYDnxS6ij/odjAZo6IhuMPj
+XILJFRILMVRgaQ5KA9TIjMubgRF/8EGn/pnjhMI9luBJQUsprY004MXM0wUbWt+SX4ajAnA147c
5EEQLdGjUArLVKMx9LRxHgJ7BZlOxaz2CedbOwA92+ftS6HaRbx7+7YSzRxRAFF1kFi+tFBRTLVg
NjYTp5aBHGXNkeSujrKAyhCYkPsktO9jpvTVeevk2UtBtyGffTssYpTCB2cAv24ZEvkZxYb/1wwy
0LUSw6gUdoMvL1nIgarXng0nrfyCED1zNHFH+DQmztNWRyTRnEVCt6rOjxkDGsIYtbQLpMJAO02+
aaHzRKDspzNWAVBgAshN5xIinx3Z2yY/R1ca0TtFKXBa4aW+69zWuFu/qR1g+eBOpoE+Z5jA/T2N
gHqfyZIN0ZkLUrMNQrXfJ+6KW83GB0phkHtgsRYZV43hhWOryvfDskcjqeSW727i/OyPrJkdstr/
QrKkC8H2lsIHM4m7MLknMVYmNVcP2CMh3L1RcGU+DlcCgJKR4l8JTzCSsD99MswIJLZG2NJQxJtI
pY7CtCzKbUf9dyhO4XDfrIJmbihJc7wyOzPssWwLiYFGIN6+DE9XEPHDD7viAcOSvwSzZ+rBOM+o
V8PO7ArFub0sa6BYaGadhb/Igueiy+BPoRabIdywlrxuu3kLYgcpVk0ZNlyBsKdseWaD2PGGXues
5onHbUtBJIbydmhL1EIjokKRr/UrVOx/drMoL3nyylau4mZGs75/GDk+Vgbt/KPH4booduEH8c6l
KYeifMnsdgBd5w7Ds+CzajjQWHlx8PYXy7QhMFQTcxgIlnRaApeC7IiffMVtmTWvuNaPHFYH+lTM
azIugj6Ke87fyaorZgC53jed5ISG+C34BJ+fChXgWSc37L3OFvkrTRKDkqC3XrKUWswxd7PPsSQT
mT09NOtJh4N6nzvF1AJJeHi5V9O/T48+YWqaEZMC+BDy43j1ePsWMkz0bpT9K972Ildy3PCiI6nY
brUTi29ZiXWj9Wb8ELob5o9r2s0aTt6kcxrYL52ljf0zvj2Xnh7Jv2V0mgGv8R/BQm9BYg8koSOU
QWhawr90EirKz/fdkEgXzglRtOSz1q3QR7PKadeqCDV7pIOF/SeDd9p5eE/cTrHbDUii8GHpJkmS
3KGdMd+nyFJ97tlCLV8uWJrIaZahE0LeMeV8Z5TfPCelExcTfIWU2MB6yQC7m4ESO8OJkITjDW8D
ciCAP2pbJLUWrwRmWr+TiszbsW86FVpid/0VpXZ9Y5C5/TBX6LYQWnFoEUNwW74I7WK1pVraKsVk
tYzd0Ac3qNcdQq67tQQfaiHpUiDmfI+/7JOaKMDJ4GiSSjFV4LeM0jocpJ1KRbtzuKbCxUaj3Xsw
RuK7SKxUaFBnQ30XHSptwgYw6MAbdQKovpQrZhOaXrc6odeAmcwGvtjPjdnFgEJU+fZp/3FLGf5C
z+RRwsDGxscThx45cN192EaR9fu81ArQWxqkFr1b9+2MV70fEFR2r9e6+hqf/eGWCjKjA8lNysKT
jeQXAkBuurQ+Gwp+pqsHCfkVlNyVFPDTUiqF5utU71frNuw4/AWb3TXeoj0tiPwz0iucRUzl3G1r
bOziIZd9ERIY57O1OTZWOVT7OYD4/HkLS2s4P4Q0UFJWXwUoStQmouzSLnJ0UkQgRNW/hRbzri8E
b24wp/Y7qLdO1I3jcxzCgWsmWnpOwwnv4IKdbKa5sIVAX+HOX0sWLuAO81Ivp4AjMR1YMju7li/9
I5QS+puh0isUEC+3j1kiXxQ0ULY+HxICO7mHFd4zstnmhF06lsdBBqy1jlWyKze+OVfitljUzKTo
835oXfsuBXazIcRZOvP9wLkao3V6jvrdlrXnyQKwOJ+6M9e4ZV4r7deSSnqXCypXBNaGQEBVRa7s
oWfdUBDlUVeLlKpdq91h/EQ+IBQQys3UacJ+nKChtTGzjQU+ja4OWef87lHTT4LATdjDFnYy8Gs/
pSJa/tGJ28RwIrZgy0hJSnwHPOtebNEzeZfFj9IYsqjtZYuiQ3sUfGCT4OBl/tdz1tVrOzNOZo4f
7hkFyh5bqG/VpV+IdIcupI9rVilyyZTKU2bhFeb4w5Rfi77pLvU/YurtDlilePY/umVOJa1arBJL
T/kLTw4do8yS9IAAWyl9lnj86f/U8ArDP0bHVbWC+ZzKibdlYUI7ByVQ+NcbxKZz/MejQnDHjCoI
mW4pgDsq7mG3dzq5lrMmIqx+Za7XC5ZB87OqEMWENhx1wJWtsqx2twwq8qEnyWYxWnIaFTCzYuDE
kn4qcYk7EHds8S1poTOMC3KcxLml3vlA3HxamfHH4j0kW+couEGJcpYlkV2pixCZd7Vog1Utt6ne
OG6uA5prFfopB1ddM0XFfOD3Pmsvlcq/64tbMOACm7/rz0DavCQNgfbCFjpgj3ROvnKRLOXa8f6k
mAwkOTbja8TUP5/H315hyaKG/H/W352zQX63lkwR2opvAGxgNh34eexa72KVursrP5XTH7I112e6
pd1Y8Ci58cOADkojd/E39KsGcZNQHAGPW7btKC1wLwM0vJUSc/HTzYT2hFwmKhCzLb1sURhfcErZ
QqLQnJ3wk9FAmcjTm14zWrm8Nli/YahuouEvVIAuNedq700d/Ys4QfXklRtWzU73bSWPCjywLKLq
LRqUw1qrsbsI8AT5U6ku7jas7qmtcgty7pbelH3ext7sPIaSQPPIcClyNkz0Z/3FvC5vte3/OfHl
5lejdTLqJdUNRBT0ZS0gbuqypuCUhwk1j1/D3EUSXJbfYRkEpk+70H/vY6l7axdLG/0AqvANMbop
fZeQ3T8r+mttyOTxN6JWzSksoT/TvC09z7N+rL3p+oYDaZj13cNksnPZq705K/zT+12rnrMHeBBk
/j6rIvAi2N+6LozRpTNoixx+9BBgwShW6VrIpJ+vp68wGEkxWiaqIREs9tnT4oqAP7T7YX+7CJG2
csHUKc3Mq+EZWF04cE//4gPUz2epZtAYzSstxOV6ThaJodEp0AdUtg4aNGdusxBgrvdlte/Ls/TV
AlgLOt4r0ZQstPJdbcnBioE9Zlhk9hyMjdGWI38NX3YRWJAQWfv9Bd66FYmPqiwZuTkwFHTbqH4D
tPNhtLghogK4ujUD0QUAUaKf3TqRBOQMYa6rsHkiC16P5doTnKW79THpUvMzseUP1siaRY0zZBNg
t0e6ooSgMcBZi+AVwDglg4+4pIW5M8CfB2rpU6QDqyU86EtlC0QO1gJqRXoqYOoiuLz0XdtKY9wX
9U/ny1nID/zyd6SpqmVE8AFRzQEfOzggSg4cqTMMzn99BdjXvK/gQVG8r50dLIPGJfu5fm57zCRm
yk+G6Tw95ks8BkGpyqGNf3WcNVgQsOJYLz+raOEzBCYxK6DK92f12+Cl58g2TETSJWK4H4NpKjiV
TmvtNmY2ZYEfYan3k1Nd6abfTMh+MTCAIAqKpOG70bdRMNZLvC52RMHNuONl3U/oEniH3raJqOw4
37CWxI3FpZbSC/j62gmTnOVDyxXYjLWyTkl4FWpUZgIvTNi+fn1NoeFUZJal6DoJ+ha0ySrqLZcY
LusZJBm7GnLjv7q6X2WMgLCluHG2ooVajwNQ1dma8X97yqoYI/2G607tiRoV8w/Z6NXRCQaEe3ux
zPXK0g4ODRTSGlZY86v1cCuKR8o+GC5Yhz45zNvRxeWk2D12PwSbcwTdx2JHaqAr7NEcgyEdFHMS
4zMshXPTEeWIj/9a5DaLb1WtExGbcpblKHNcx2uhitE5BdfBb25iebRaN0qoYAd9LDjq0mhbiuG/
+d82t8bsaZ5cc3MfyXPElxS2R9K3tYuCtjRWE1uCtlqMFVNDXFxz5nEaA11CmVFNX+TZnEKQP1Uk
e28dWe9ijw80NFP5TN7YnJNp32XPU+tNJj7sDi9CSRYh8cX1wqtJ0uxUGSzhHTW9tHZkIIJVOQGK
ts7i3yOPm5m9rejwY2vXRd73IsH+vtuwHl2JD7AimybsmSz5G9EvAgEq3tlJwgiZhTZlscvkoImu
7k8L0IUmhe7ZCyM/fIKWh0FHswbpGVifSaIdMZxzZDlua77UWnYeQPFF/BP4lV9CSro50hv9l75U
kVlbNBuwLBqI8YO1waaffSBhzgzQ+3MRAeJJgchbvlGle3NkX0hB+pb7m46xS7WpCTkot89r0dGr
L0IWW73obZaJhc7wjWBfCYUcUDJH6+R+TGKIioRamvNz/OA7ofyKFNiJDk8jDzJMTaszaVWzLob/
hUexDFhVGghgkhyjzWPg7BQrUgOm4y+px/ttxwxsZaI3BRjZM6exYl5oI0vyjyMHx2pRmuF/LuWq
jt5kezrCn6Tx6Q0s30C57sfGpLIg51mC128PwOKxzhJbCQba8aiJ5WqSlr3YwlyaEvLDhxWrGHS5
EGjmFQCiSOY/E2jYShngY868VBy1Th3PLwGRuq65nSvvmm4SAB3vPaicd83CLK/8hm82JODiUkzS
6zh5T+d0Hh+57I7ErKyNhKWqpikNdpj+m5+q8t0JryPmyDuUuQ8zRpt3qZR1Wry0FOAX0nInzWoM
FNYHfMWtdZ7V634JtHl2P4RjPtR4nIpf+p02HeclFFIB2EwfRWmWsm2INtH5c1eba6vyKDe+jrJ1
Nvc3aElFSQTcGLHp98IjpOOQZ7+DF+G+GUSOJUg6T4igO22SAV0giaI3Rvj1i1CBoKdfB4ARE5DP
sIskTRTTsMd5Kc+yElHGy+lkJdlh6I09tLg9M/aSCedthqKlhL8saAfymrRxwOnThF26V084bhpv
/mvr6+6drt6b34dVLybXiPkybUhgC1QZX63UIa0KnYwrlbMidf1NitbOtcpcPuRNJWYbVBzR9wTZ
0hjk6wtmtaJpRTy3DzpssbmMAhEL0SjZIaJ3+9tYV2lTy7yf9alp2b+Zu7dXzm82Iooas5L+HdWd
LSi9kCxSjJY84Jtv0ituwpaaeF609f9uisIPaZupwTsEFcD5jJwOIc30Hps2FxPko8UR1FzSa/36
XqPqVrfwXTUb8w0C3hGpcnCxwhkRnEvtGXb/tJhX4KCPmWR7Ztb1RBzbPe+wBHQg5wxxw7xbMX6e
dBtlKoI8OpyqvjL9mSZosN2VZclpmdblkXZ+/jCnVKb31OHqGXuIBmF5gy2Z4QDMhv7EHpHaTsO+
CbEzqmbavBnFE1/WEUvtSIR8NrJV9+0Q5n+1IHhIHweNwSwC6IbgacRiLARYYQH/9iGX7fQ3hmGC
RfGYNHqnnp54usnj8PIboxY2hnNzbaF6UNidyVaQw3xxi0EEqZHMe/bkxbUNfZcMy2atwrsTcgSm
v4dlucdoLckiLL1YRoF7mb5uKq/UJ7XGodQpbRUSzMMJP8Vhq630NC6s+JsHb/idJj3OEF5+7M0G
GnhU5aDIWODVzKPSwrnS5XOKzF3gsDrCaxbIYHMfMCfDGEzgv7ZJApXf1T5FY2SG5yW9w74upswe
eGdyKosXcUxbX8ZsUpunspKv/HtgbFREjGz1xs0NOWafDb608qh1Sdhojsyg8cqdbR3MzkGV1AWp
lN1Bh+/rac2CGYxvEp/V8yQNYRoGrVWM45sGvlLJ59pJRSfRG9gETRcRaF5QU9E9Bkd9lig3vhSg
A1IXefOckz2cJg/o0+zFomm0VpGRKw1517cJMQ6cO2JttdwfAgT4KWHLLsNTYkQnShJXl0C+kDhO
JEz57VrnkF0HaAdOr4x2efKWVEDcE0mvU35698kjjgRFm3HEpm6KJ8+q4VFcd1szFY0O3Gu8nMHi
vQa6VyTnrISNAzuUo/gcOIdlXfTSRNp8EpyhraPSR6jXtwBoEL0K5Cfo/Ts/dCVMcjvo8ALvXb33
tlLOIMm4QP7uUKOP8/4rURcQdYfMLkUEaeyuFpunyQzUD+NMS7dW3nJK7dEq/QA5jN6UbibS1qZA
gNR2yBxH7YEHFhjIbTD0uA6KDVSbqkXjlJrfXNCkMi7z3UhC0xOreT5xmu7GKeMNuGo9JWUdMVtS
XEQyvLHBv6wPT0bEASAQbBEX+1McJdSCwlijZ3PTlF68IAUbSWterq/+U9zBvTzNdazWExH1uSek
30DL4mzRI5JrVOlz1gUAjRKmxChadtDo2t0CuIiq8qurMBuy7etVqzK+b3BVgel2YJYaBPlOmlvZ
SCy0C4Cy1RVIpqrZxv8DgCYXEfg1ogGSWqe4x2oNWqP4O6nvzNk63rgxsTFx0auPNzUjvRz2nSQ5
VRPn78ZzuGcQ228xeb+Ifp4xz6/zfv26l+uMZxbgXG6cyZ9X3uFDVq4qH1MWBKSx/1gs20IO2OFB
3TLoRPusH4ZafUX03uw8S/VEpzuaCHZNabSx89q3CEcktbKegR40O8MQ1HIb2ID6mVTIHiVGLFCn
1Nm0eK5yfkr4DJVa09ZQBrrz3gksnbrdqXU7ShhYIWxuQwY0bsBeISHLKQIMZ8QQXV/Gv6jl9N9y
DZvFKoKbto++DkpuHQSgdI2IHelwzyog86wKNs82mFvmG5+9sv4AZRUUL90xgPtM33hLKt/52mFZ
Pa2VKzs1NaE47jPQPGke8Omnt02j9HzK+LQFoS4xFIwwF2t7hMcXTumlDtDukFvp3HZjDo61AFTK
EHC4UuDgp7btKgrLrIOFhFCMLCzemH/DkmvLK6l4/461oDgh7cPKbHry7hE1TrcABOevqX6Ugn8T
N6rMsR7bxV6Z4OEWoT8v/OC6f5QCVUwKsEHRhj+8Rc2k5nKLVF/VZAdGyPHiXn1Ed7cI/u45X6CO
8uPt7BrcKU2wARHcJFox2WaXkJ4ML1PquQcfh86r7WFsN0YDDrJCwiexDJ+gUepLE/cWhWOCmd48
PF1HMgr7AA4Nm5sWj60AH6f7AIKUMOm3grva3SzXoqBDfRXPlvEEvnIKeOd5qewYd08SkftbGvyd
gtNK0sMjXVkMXRDd0aUiMXoYYcfcQbgSkcaYzttByFP2GgfQXXlDlfkM4HXPLeJ/zji1NNX50oFR
Sr67ddM6axpSmYIlcNVNFgpCXqebll8gZI+qmgLD8CMR0BX7OE5iUnpV0JGxBmDBPbE/dGcLf75q
a2vfBswYgVT5saFX5ZRc1JbFHcK1ywj/24Cy4VcQPUw8Nt5ZJ2qrEi1ZrTkk915dcdFwbawJUZTG
fjmrk1K0puv9+tP/5r+WvIw+ynmMV2oyWk5W4/T2ymHZj8EIhGQkxI31DMMaAUpo56iqMsOwiCtU
e1tILe09p+qdRgBPcWEEGk5ZkKbpAENgWDIvcub5okLl5ghAM9xYEi25AQ6f1uQBEt6WBVKjwmxh
xYXaCoGHnb1u4KevtjRFUsSDXrQXi2lSzojIfm8WICSpSp6h/dgSst6QzStUtFq3BLrCPNvSDGfU
JxFkOQs2irQm1DuAVn1O182exv0SHB0W4XHzT61cXiIIsRV3XrojTuSeCKltdr0QoVo08spkD56n
6CkIAl9UJWuaTttABSp/ZhKLTTL5afv/uvT2Qrt+SM4SaQ1j0b0jNiHgcVaVMMz7VNXldWL4nO71
ihoHh5RhysvclUWpTw2J/zN4PxNw8t03FES1I4Fsb/X6/R17A57gy2S+GUp4W/xbU3JIYd/e4Hag
xGXaArDpblA6g6gUEhu3v2GA7d75J8kvp1uafF8IVWqi6RHkSsjYF2yozqvdwcA4lC1EFfW0oBC2
ZYh8momV+lKs8kI/ABVkHIy4pvoGMU6U5sGpu7D8rif0o5NfrKzqSk9DyhCmagc1SdznD3z4hW0o
L98CeTYIJYAWT+5QJi6UTBXrCvnIgm0RRBSxOd34t807iq62PZaQ0ZyN8pZDt84vOiVh4P+FTOTy
Vgq0YPgmsZtEcaVGUQUP+QQco26imEfgs7CDd+cm7awXJCAUvetoqUPb01ZO56Zzme5SW7vJhb/G
v30f6+CZeD4vbH9ZVpjS49+mwL3BUUjKA7fO5uxETv0H5UXSKI/lYUw9bj9E3UVZk5q/GnWMC6dL
z2ken6Cc2f0JwhnRDjwBb7inN4r358CaTx9UQZajD7hyfNZDWOCtq0HlaXx688LwmPxVvWLbP1r+
agWtNy9v5EkoIQE9HYDG7fSP18MeRQ2tUs10HVKtzMqesfVsOWik/IWK6tPayH8AAX/++n2o9Gba
25PsnJX7jOYkWfkGVFaK12dj9E5lrwHwFlunQDrkBorKWbCg1A15wR9SexI9/gGRrn2bqPon+EtM
N7YYbr06E71TVrJZBuM5U2JJ+1ewdgL3h+2gZEua3PBjk8jPECj/ZtYNFmOOiCA64Kotu1KdWXqf
xXvIm3Okfeu6CTvNxO3nSSJPImmyPcta7GnTGwaBcErDmD/xfFJcbX98TrFg18rV+b09hCBdPnFw
WTTTxaSYG9oYIWT/8TF3W4Fs4s2wPpMYbNL/2XDpQGY/g6H5X+2a2nLRnxn0FcjCymWvUzQBVt4m
QP2r+3stSnoW1RNIHAVY2rAUx0inyX07jc+KZdiYb/s+aX+eHzqE/i/j2Ix22oUCvAi2OtYCTSZU
tkrsPjSt64nYSVGyD07wXu2gsq/a8XFyH/DR5O1dQLDUm9WhzUUSYMp/STJ8tF11Gg8IwoOQyuDM
PLRndLEXxGaJEVgpXy5SSvXZ0/Y82xUMgi5eenkfPnQqe2QdffhhLmQkzuWLgCPu07f9BkIQ755H
pPtpK6hL9iwL3dk22GT8KV2DmHnFoGkWMLCoPrmc3480NXni+DNlse86YEFaVIhsASYClVvr6OoK
GzKIey9JuyxfiucSyPj6odAtq+eOVT8NNGgKj5nSfykCwvDsSqKPksJjSJV9VN6pfYJpvL4sjf5o
QIKpQUxFjJ55nkL9g5UC6Etieet1EsQpb+eG3k7lSU5rnqnJ7nLbLUyYugrWHv8tSoQwD9puwkSf
RzE5UCbrPxGSAv4NI8uUg/Tlb2vK0kHyijBycTvlF/ta+3Zknv5wVoLX4f9L3sqGTFhG86DWzmdi
x7Ipunn414RmICFqf1HzVw3hYWTwoj7PrSIBma2PIyqZx75oRoszJ7IyRjm8HJRL8ds6cz0gqTmU
mYFKHM5/Hd3+pdvLzTSCHprl6RsmAWUDQAOQ7Mv9CBJNbxBGcpvCvlADn7OVcrGimku0usk2/K2+
nHdEb/sAqxk/6aAiXTbr7FksiUqeMgOMTLHrXK6DpZKbhCRYQn+d1GSpWKbo82O5upFVDKgSTpQz
6+6Q0EsxbeIjOxxzI8KKFlSHC2M4mObLfMaDA3iFsZOHJrkD8D+ssuozFX7H7jHnzU1nI8sr2IZk
nIro3bC5pf6znY7mjwM+4el6J36npJp/9IBFNyvlSdUxhn9SOYAcByKVGXGMyvgU5qZIi+ArAf67
qJqETcpUjONRF7aC4Lwn7YmM9KqhybJftwS4FUR2FwgJct55S4c8NlfBYPPiA/FMkqFYxy2Ow3x9
pfwrrA5pzWs8mlhYGg7pHG+xkdfA8vT8Xaj9zFRGKGyeT6lVm64f/KBEU/3ECk9GpTytxjAiO2lz
Dov50gruSwo3WjcDVk/A0WO9UXlH41J7D1Yj2Zr7kszLqIH12EAXi40tx/M8OrEfdvLcjEvp6man
zoPCJCE5I2649zM7UgqhE1y9cWlxrOYwJtI4Bb3iyrHuiAzt9812BimrZdtU8BHThjW39HBfej+O
PKrCiA8LRR399RD4LfJItLPoSF/NuWKnTniBLTnMdr5YG0iC66nS4qlmOW9r6tAMQIMVN7lkhe+d
UkT7/SrwY/jEJQ9W64wxIOnmvqAjd7yMQ8gRAu6SKHDAKgkLQYO2/5dAgzk/ZzjZgCn3xN507xlm
pLXOp3EksrUiJWLDXH21IrW+cs3mIoP8lfgQHrQc+D+tELGCRK6IU1efW296xfsunCGBKQwEiGWY
nm0x0QSukL3muk28pA+P8GMkjSYJ0CAuBTwWFvmuGKVnaCIgAGSObFOdB39ruQJcXLwjJrFRNjM8
DSsfZi2KlgDEurVOMQ4Md+YSMpJ1dzZTJl1hRGQeJnbI3GE8bVqSvBY5a6SlKRfBPm+n7kgad0Q3
Dbue3oEAx4WRrjXka6pgROxBdpdSf1CMltfSSA/GC6hc7u2Dw39Yh1oBTvTe/oKhnp9KjZXAk4iK
tALxf4RS3J7lIdr9XLrBwbUlEdI2yiM/fgpkFPSsxSAmH86w+l0ClZTQia+lKYMvDvVX4PSkMyKG
txONyef/JUoWrCO/+O3IGIXqv6U9xOkymXVPhoYwjxy0XM+/pe3Czc59XUJCiw8C7G8FrbmEXbKm
7SqaLHsaM9k5PYAxmEY5dYqfrgzxBFVE6AoAgHrcct/k+G9OLC1DX9Km90/bh1FzbytQQ37vWr+y
j0BsXfoHA8qZHu/cbHgqdd2wTVsFNh0jrAqoyn8v8/wGar6xuVMy9ZXXM9H+FwxZbk7GNT0hH2V5
ll9ssHw613Lc+bkhOWnr2nqVj+MztwR1WOLNaCzXQuufMH/I/Vm848wZfKthhUcoDIaBYzjyRFEN
dRDFEXUQHxk1cuCOzEk1ADYf2u/YZ+x3rXqzFxOWC815ZJJJtNDJQ+cNVfR8vs0n2aC9HyojrbI9
IsYXNSKHRxGvlLQ3GDfcR3bTijEoNvEBg6k9KC4iLlda8MFzgiqMv2NB6quoInr6mF19oO/Bxq4s
q4Efd0lCGIlXCaufxspS47aBkg9PBy4J42LVZeGP9P80EbfqiPUsqnYWnkpZ8/nTBsBlDR/2Nfiz
SkXYwZjQcwqhd+Po9E0UI6eNFgr5eqerbmq95WVm3v07lcY8mp1+9B5jCi7EYrzXGV8ntHn/6wfq
A94GSOzNi3iTmn2RWUFBg3mccJqQ/0AsyEDYAEw4/SelrH19rQ/ZFQr46Sb/FV0mwbiTdrZuIj5E
m2rcGR/AriEj8P9C/C6QuRO60f+tRsacwoK+4m0fpdl7ZJUnLnyhb5TxCzGthFX9AqWEnaTmaMWI
twuMF2qxTJMZycUb+I3wsBjJt+z4MGea9k51uKlZ9k1ae3/HzcsrWqQHasnRSBnF9NZtQFa8Zqbw
AtRjYnwbYz+zzC60uanDpcE2ty93XQk8lF+tXpGp4GKYcHuw+asm54alU10qvYZWBE4jw1eZWRDe
HiF5bjm+lUazKjJxUIPZC6RcO/vKzPZCHnqUz+VbTpSdzVd7bKyjWitrNZ0/froqWYXGjBkP3jVr
z9g5x0msflV0n1QQNAgyd+R4ZijBGuRYRmk+EHAeXbv1CKIpuxsC5sNjREOa788smyzeADhbJH0C
PxjftaoPxEN0/kbOzUK95422V/XgYMXZJHPcMal1R4gl/IZX/hm2FDHPwcG0SU95UlF9OtzCNTxA
rJT7whagLL/P5cUR6aZAMjzBEbTaB6quCQ/Is7q4BltMivjJkWNzq8OpyCkVDambtEQnJkrqm0Qv
/w5yl/oiPOP2bYM/xETKvE8Z//33tIfj5NuyqtnZCmY+KOqQVRKRBZOryz6BMaL8piV2uIOm8LH3
/+HQnrWFy+yoHXAIHwBtd7UGIv6y4gf8Cxrs3ifGkeP/XTS/sbuPyEFSOi4HMp2vbnfkkI7YwXKr
YDKAWbjXPBBfz/Z5ykI0l0MtlWVDqRHNnO3CRdDq9PFS7cJB9DTBqehaX6vc324Kz++M2cT0RJ5+
9jdAUyjNVGLkTT3qCfuOk3JyIsYdPyUXJKXil/zXL9PpQ4K2qlIoa0YoX43JQVuz0lRO8bd3gVPL
Exr16x/iwtkm+G8az9NJHaJYpIREFxMB7FXBuaPFyr1ILmaMs2MloZSPR71o9YbqlLGj9DUcCktU
aK6XewyNA4b7Jau9FIPduoHz7caSzRKX1VAB851iN7yR34X+3R0ujuaFRvkGg0Omr6bbA66qH6FW
qhj6wS+6zXwk6NbMsz/AXJPxC6ruPVnIPoIUwdTPw2o8Y0KBbsl9mhOTM1s9oZFLW2VMVfqCEkWU
fs+Ti2MKt60h3V+qZYkN7C7/edcU3xXx8LR2YUzwADuubgy4K//FS3yfc36UDIdRc8cw6R+Zrg+u
PXXubm9f98tJHrsHTAfnAPSpGFoGyoTAqqzkdzfHsJC2883u/KMT5d2vqk9zHcu/HrG8ONSaYZqV
ZdH8RYQ6fLWBGoIxRefgkV8zTJBQyF9ywK87Jhr8NBVkR6tM76hQk6ZUYjrO2mmGQJXJKRJIonz6
JMhykjfs0vMWqAtOZDAD5LA6QBba3T4WcMbLTOr0p9U3zqfBistNomAITKIYGsPi1EXdIoa7gGeC
F79aD5kpcovrQCT0Yfo5TIqfXGNBu0D6iYpAXAWzjsTcAGgDKJw9nsYu4iFjZ1qiZ+yrNnB9rWXl
DSsqYHwos4HlxUFwrauDWhNv10BSCGG4t90MxgDP2N19Ywxe2FGymh/igR8B3NXeT8pF4aTH8Z5s
8ZiSw+DPoMGO9yBEghE+E21HllsLtSYzlZcyk9fSp4B56yIacXMnjHTsXTW2RJ6mZU/rv0v8XXHF
FkW4+sDsAnmuI56rEIbYA45L0MwAeaJC+hmpjRp/AUFRlnp7PUMNn2MUEAu9X8dtaf/27D3mixea
yfU9Nfa4swNOej3ED/Y2z5UB79tImBGVd2dA4A5ZJoM6KpYklwlGKh2l6dcXTDdhYcChm1zRBMP3
bC5jweRaLmiltm/MpzcN+qa17rhYb9rHZq1wnzb0/Hqg5aXH6sWPgXOXEp6vXS8u+1NDKQck5XZh
Yuw6G6ohDKpHTEaV70nsHQ5NLCd33NYGVViMvSLnalQ4R7wL3qQGIhkuBG8e6hF1D7DTRuybTXeB
KqNmlyOipkv5kbm020oigNfz7DwntCQ8+3KlUn7UHKuOsH2e0NqWmrdv9pNdmI49zKklJ87XfSQb
1W4rKHkmDM2OglYpxDb1iZouEa4aCJvmNAte+9orR690TwsxFlRHWEY5XpyTyn9TUpo97G7IDxOX
EW88KAdQvjP8iuQk/X6WOIm1uXi0lbCd+IsFsztAHaR2lIxbQASNXPVylj4JeT6DGR9BlQQ3p9af
Gbe0ZlPaUBgft3L4EmI3zccOtMjenXLcG8yd48emSfD36OAvI4F0d9S0auq3Q4PZU1CEx6sH0B2P
rWhy0q+cKv9Zbfdufx7QXVub1Z04BlWD3aQg+K+h/I1WnmqwYT0xzt5qv9Dki9TD+dqJVncjfKV2
lEjjT7Hu8u3pRY6wEBD8cmgEEYu3Nx3CwHVNM3GGHblkaLT1KllqONLLyitWj5EtTW0hYsPMHobT
A0MDuqb0NdbGg7sS43MvpovGydRmY7ZEjuexnMcgI3WDPh0P81/3PHa/47bFZT8WSQxoq0FN9g2h
7uu01QL+0yXoIIHRJi3qPaY+cAfu6JcAxvYRkQzxbSsSjvIs98OwwpDofHHwPT/OZFvg0coqMuL8
FbA0crnMavL5PAwcXsb9AwR6gX/fa6IymLl3wTwdaOGqQLLYNFA0uMgPI0TgUfFZ4JEg1BSH8N64
C5NOrjtl5Q6vfU+oq09tG0Tk04NhuoK8lkKUF4JmQUWJ8BtCC9cOdP8QGdK3wRWOwlQrvzHG9A1T
jc3JbqpEIrB5dFALbbmjU4OrmckMH+ZKQhVbZNCKOHYaS80CdmT7dL5Sct3eQi8wb4sC1y03XqM3
13JFPwkCj2mWi8QfEGkNHqWisFwT88wp8xJUxrKpfacR+NGP0jc8mhr3xw4ER5NmU8j0SQjJqQhu
xrW+5R4fIGqm+yrajS2LFD5ncs2EzYD1Yw7jn7oKuNs7zUr1leyLrOCFIZdzryIIzckLMIZTepLC
PX2Ug5JV6f3paMvBrq2TgsJYSjnCu3H1jrQsUOSqmimckKZq4dnADwhBJxbK9k4LGlMsPfQvgxGj
F05Jk6mNQG9HyE2aVVgIzRDhWkkDYlshvYZb5xPAqXSi3PU6lfwZVE9WOU0SupeBz89TpeaeVboK
aToK2dKyEkgHzjsQjn14MOGWjhCjfupJTEixo3TohHH5EEw9APe3uSoBYEO5piFDZYO+qvA7Exp5
L5ZTSNGz/gfkbYl8qusrH20s+blr5zAKBXc+s4etJYZ3LgmsuSB1B3N9zUSQaxaYv1pWS9BfNjZS
RwJcbqu+p1qDB6a6Qv0rAdSh1CSiVXAu6qQ39LfQmUT2zgH8Nik0HD6JOBFPlDt0DhL7fgI6Fh8s
yCRQcRnLq05NoVTA/dJkpfeVkGDTYFkFm5mkedf9vN5mdK/wUjNfjsCRsiTLO8iFN5o8TOYz/6u9
Ruhb5wCOrU4/iLTwf4cOQ+1S7TUm/a5f3OOn1b6ts/UscSAgq62lV27GvJXqEs+fL5zeN/MsPF7g
gy4tofwpsDxy/Pn3lx1l2bQN/+uvs4ZRQg26ixFXOMsWM4D/40H5Efb/c3mRjxo40i82x/4kOvEE
8Ut/9REIrCgIMIbEXtKiX/+RpXgBW6WMuSBs9eYhYRwibdSndZkU5UR3iiaHSN5u//gKCKmHPWO4
nJeHcJti8p4EQndUYeldOFZ6ThL1N9jjOJWi5x6kkI6Yhi1Pa2hjXkNeJiwEs7XfPstplJKqkNN0
HU2EaHxlezHD7knIj9U5RQWmYetRcGeSkd5pMRqbc8cX8umDOAiPeXkgCGqgjkMMFYJGrIgsM85o
wJu/maJo4/PJHtC0kPzPrl4wBFBbPGa5A0pUGpSpjApvZyMw6yuBYRYhenaamEmW/eZMVunG8Nvw
oIh4FB42Z/Vt2DuJnYG2vYpc0wlHzt4mlGpeR/67OQF+iXZDDOUByTLq4kqypETusF2CHH5GmYg0
Qaj3v/FwsZ2Rm2X1+loFt4X8LTD1M/5+cLs3fEzeS6es9jvDhEqdcNL4NT0RzQ4mSrtUnrBfG1D/
aaoLY9cI/ifL0KC6WZEdpUCIkNy1XQrLJ42gZNKMb+91hK7+ywlwdP63tyTtd4WRk1gTRcOhRQV8
ueMT8tFce+zYxI8buXdXP0LGyR3dxVNygy0b9xtEMt001nVHA3f9NXNuVYVLYN3sAh7Zg5rY3xi6
xbl1VgQXb0JJAfbWsm3MkB6HRyhBoLg7PXHbzPr78ZnLEImmYviFAMdB0WvYHJe+g8XC1L+U6mPu
a1cr8nMeC5f7Q3XpFvXIv8kSVOrfjrPlaDOS+k/oNJWfyMil0HxwcdimUWV0/kwqEyqr5jETgypY
XzzZfn9qTMP3wS50Gy+S1R1rA+3uI8NCapOkf1kWoBOVG9wK6insMsiP6Z5IJC3Iin9wwfMS9jra
RULEqoeJ1cFtIwTViXIfaeiUZ7bmmDl5YBDd/PVafYesX/xPWp5h4CzBfzmshXC5SyqHYG1OkKUY
XrDgyeTFTJpOfBvGlbk0uMvJp1zy/9ox24xv3QM7IX9S3HsZDrXKEmXIhcCdxB08yCTNt7ZDoiJi
fdd0yjDbDiVS+NtXqUj8YBvlcS7qANoalj/TcUNj7IodCh6Ou0poc1oE/5kY0gkntnzOiUgok5j7
SRAbHCCZdkOuuDzwFWKwmviTF9mqw5AXwjn939f6ANSb8hHALF4AEP7BDQVZPLmtuSfieXOnSCr7
fnFLznVXpiTPBxylKFk1Gn+4Rj1YUtIJXmqX1ZCssHBxxF4nepurW0yL3XnWIJj9QvfQdX30/l7v
xvsvffh5oj3bQhDCwhscxilSFs9+SBteoLv7V5yGhr8fLlAhCo8MoaEjtPUwPLc98md11LzotEiE
61xV62Fw+xTOm2Kj0doYI7B+OzcFwemuSSuBn4z+Ix6PJo5ibI7K4KEqDrjWyMlzQQishWHrtlxK
S9dVq6I8bTlCAdh5G/jQx15ruCOYEVtUuFlPnjZ3qXhgK2NoTCMeN0P97xJ6qiJESi2YF67ps1Ca
QZHaHO2jPkJ5YxvWuUQyIleA3VYSnJ30iEw1pZQEGjmyLE6Ny+nSUlsgGpeOwZDQfeHXUvco0Ee7
k9KdASQjjMhTKd4Y1w6bm1mpCFZ7Pik8DybTFrvRPEmtDliNOA8Qae+2QeME7tmDzskgXXc1DJXV
bCt4jVA8Qkvd8xnvJ0RAtRduw0f8N9ROe1LYmiizbFYIySmyCpI8VDOpjKJFS+N9C+PNNmvcpBRZ
mUU/FLln7vg+1kQAqOhXwX5FDqcZhld0eovzHUORgCJ8DwJt1YTaDGDUDanoPcmTIQiBwsI8iEtA
t/iWJn0tiOdiPaJ5XwPVRSz0XXqNQ/piV3m35umtGS0wfQcY3EmZMIgomCuAPtZFpnmLkF8YwwTd
QeR8runA46QWoFe8vWdYAOAiDQJQ1rtFMjkbkJVFfmC6TVq7Z44nZepmoPgWbf/HVZ6AOUJ7nRx6
xXrg6jHp20/eCnSNy7CYXvWq3onwpA8WBnfN2Ia/BdVfV9jCLqWonxcfp+J1gFXndFzhaaDpeNjk
jXYd6JQOi4RO2gT93pap4L0+E57ceMw1z2gcQ5ycAIiHaKaTkYXe+yFmj8fbFXEE7iJbEC3cC7xI
SQlGwanPH8K6UIrPQl7g6p9mq8c4j+fQ6wR24LiqQ8Gaz7mawm2hGB8A3Hli5/OeZD3LwE24JDvA
i5vM4YjuRj3481Wn6RZRB02AGniUvqyQXxATaZR7pOveRTm6TN0mPJ0tSUt/G6oRCQwCg8UBPMOo
g97bm/EcxQlEg8xJmJwA+Nx6NsbYhfdaNSVp/AiLmdGOnZFL0shV9nEJxal+Ua2hVpvhs/KgLPw/
LOQAI+RmaV244lm/9vf29LqH/bc5Qw8vp/l7bT37LUEQilY9viyp2RcmwXwGt6WdtSNaFCkSih1a
cMRBLOlokAb9tdhuy7o9kqo7mLrsd9NCPn+MLXN2rrfAlfwd3lUX53UzpaAiYKC/U1HDRgm8cx4Y
ps2dmReA8rjmsoAsZw+Ze+iCOvaV6rJl2UU4SbH/0S7YIHqD0xNNiMQRqOxo9OHXBv+gF8YGkMQU
wsMMdCjBqnypGOT8mOmlg7NDtAzxh5m1d5O7L7sUDzjJscBCg8PuxORbEDF37bAazsK7iEEsRymn
vZB08Mv8CfRI9DQlDVkdEm6AVICX7PcpPUiN8IkjN4GkXcFpgc+qG+dMWGtFkwu+JjVYYRig+V39
ynjNhqiUgx3zBrV50d9f+htJ+6FB2LJIueNG7WeCv04/C9ZihTK0ETeKWQuhkm2olhrORPoADY+U
WMbq+3U6FAWyvepuVsqkMy07q6DggX6sv67cRDAbfIDmFMgxjdD1N5KZC51c9YoSLNaa+kaomUvN
3dKS7ko1n8K8b/SYIIor7HFg993sjxrrN4PpT2fXQNpmnsHC4ODq9nBgxskCrsXIaI/A2GFU3Uel
CUF+4YNVIKo0Crj+nedYA1L5IfE/2TMxkecDhQvOGfDbSfkoJNZBWleL0cvc88DmLsVc+MXwAAqN
ga2rc+uFbN6XSwe2lKULlNjayCi8LAW4Tb6MZ10MAbgREf9KLsjrUFl26KbCbXP7p+1oane0faXQ
p8ADkRlb/onTF4aNXWE+ST1VaLRyB+TTFY2ctwN3a7oaBjCiSWgKKqoivmjftRVhlGmoWYkZB211
hvF1G1gL/8Ag6tE2BRyD3b0KEvgmRF+NKoyrJE2D5vdOg/hRI/kQFI7Smskk7sQv6QKTtKL0lACO
WJvKgL5aus866YqRUimN57TO74VC+Z1M7oka3tZXMTMbBG1OfAUYgQ+kZE+7iXiTgi9lqtmuRSEx
+rFPdzo0JLWShSuMx4g+6TnPh8oONwEkMza9UZa8mj/pXdJ+RUYFVZg29TTOurM3UUlek7Q4qAZ4
mpSK8+pdvXELRJrd9RJq78CvWxUxe44AW+ZPgmMlz2YJq9BxM6gcPVtQ728xlDy97BQsgutH6gOx
/BcEq4r3LUQVycNEFEB/wOu9LllmbmFWg2qMoZKD5jWqlNXSVAOkyg5mwRGBAndmzurlqOfbv+CZ
8BYgFPO7k4b4XLvZWg1jpQ2JU4IAJ01KqeWbr5t7LM3DBRUdvorNrnteRm+TDxDx08bFWc9FdFqT
I7MWTvkOezPYvEsqlZMNvXqYrYXogwAqL87ZAgStGdWYeVbr1TlPD57XFGKHpZlckjpi4kvjV2x3
bRt0BFOLznwQeJ9IkovjT5xtgR+IsB+OEGyH0Wfp2nLKxzHGxDRskYzvircBRXfoa6lpd96oQIz7
fekK/bJ7f04n/Rn/OpsSqXYJ3kXJqoY0jl2TWmgf8MJQms4+S1yKxyo5ZfUPP6oduyZznY/XD7tw
Y90SlFEflDyDl4H/6QGTRQggAdpw2UVTL3JzUfBHR7yvlp5KycfQY9JjCbDiTD0ngszKgyl1zUIV
USDXcYgrvyi0mOsgwgAUBDj9XYVM4/J5/Us31S8Lq/a8uWvCe5lrl4l9KiwN21o32McsG5//LvKp
43AwJy/ri9xueIM77SZnDuTRSHh5SpL80QEzDBqT0iDAvzLpj+PTqX/qWv8wOuRUUf9CjyXZeQm3
8Qc9EWhwmuL9yIdVsseIpB7B0l+QmKrauTYN5NbLEvMWMPY+D8+2CxpYQ+yfKeikjEPxLSmCM1P2
8hTpeqT1RGystAABvHkOk5zNaH9RNnKaPRIl4JwW32RhHuU2DjV++BEy7vA7ZCU7XratJLAtZ1nn
TUheD/3grM6lHfjPAwfJMBTyj4O1JZh0IZlsM3mDCH+R0HVratN7okVDgHiLabFbiGSXnTZszjPs
ihmz/+84MTEHF4O806LRa4monFJHJYU+osVMm8bCdrp5DKjye382rQXtCmH3aSZbl0UykcgyYm/F
si/YI+XFntpjDXKUYE6vVUTa1EP0hgGeB//83p/cOpeF5jUHYEVgUR+SqT4pEeIqNI7TorM3UkdV
buci4lu3/LEpeBW3DeoIIIhFl3p5eTZewg+spto0tzbfMZr1paZfkpz/o8O3x23A+DTIDrL5jKdk
xyrAbaDB2gRp46D4uuJx2CJmexQ2x+f3cs1kVZD9BVmWVp7x1CtYi0GZhOFzVZBXTHmtswc/9evd
iKNTrNxbsSFHU+JJ7jDIKEVxnVoHQK9/DafpAPNWy6HKiK4uUSD7emwnxi1ooA/PRhaEchzNufRO
+Qlccnl9cUZk9mkNiR9e9u8OzRzcGmkWo+bXU/lo/IF1e+HUaF3AKh4S/uVKrkung+ashGURYsfu
1RE3/RFtyx+qLID3ZaXAB9MC1a+KVGP2da7uL0XDffUsZhX/DHjxIzg5ET08Pb2kx2sN+lUicyOa
dftUlKC37c8ULaxuZmb3sCl4g55CUQaWRw10Vb6Mo7vq7ALH5A/UnNEDk+GmR/rZ2hlVBrv/uKRN
P8ehOhc1TdEGLxGUC2PIlmXPj5ZRjPX3HhpLqmMBl8BOU3wXlHZx1QQPhoGEsGXzcl16mD7MoZsL
ydcldNJ7jTM0yBjLbQEVMFVvJTkTP1DbaEtc0or558mrrsXAu+8WxdhR6LZprEdsOA7+UEvC3Irt
o+uFHJnxko0rOT0zMXEOicbT5JuNLuwcAM/pBXpiB+/2izLHA02tI+X6+S0vobmGwyROgmtHo9Ha
/7GQb7xggqXL27Cdm+/EmO4ggz4ADUyCfqdeNa830BkRxDLC7aoBDaGV0afHr5T4nU6yGu71WSjT
ZTH3P5fT1c6X8tVWZrWwmLalJGeun7Ae9054qF1r8OoiLlvraXDMCJI4a+jUz5ksF73jGuMw4wx+
8FrNQR5a99xo71uiRrrkOY2+apEzu1QKhCsoDiYmQKblwjSOKiLc6vuOo/aFSLcquwL6A6F8Ulfu
5GWpgDeV/mfJgiHd3A/wzmiUXYsLFouT2cA93gQfL+EVmvsQxIy2D5MKqIDCV/wAGL4036GhuYk9
btCFe1d5Z2/vqw7LannFZV3cw2iuJWNTz3j6Ilo+onQq5/CIbjHFHcK9CdfEpEAK2vv9ohhCA6bs
RG69eaBkJwKoP2UrliWt6YbgKrqKG3YwxXtflsKh+PkytXtYjKZESzhOuAXOIfBgPHrksoraTLkN
4LHpscOcGMMcBYzT3undNQKanw/+hB9XEh1foIj7YbwnhZUpSXNZCkeXOFSflfysmGHJ25TRn0Zi
YO2pNJU009RBPs8A0aZ6cU52l0fLt5f+zQ5OtrWd3lpAN2lxCMgbkX2CbTW1DOWyyo2IoblBG6lS
tRnUbP238a9yhP5cRd/q1MNkEikaSWIusBp/+hSe1NeCJWmNvAcNjHMttX50vj68myJMJI0KzinH
yCL7I55WsCyFI0a2rgiMY+BqgURlDKqonm6tujmQtovU6hsn2TuYX4HNBweAnTGFhiRyz04nTSPM
Pa8Ifb400X51HvRZ+XRagz7sqLPVfcl3A6NdZKjcrpx/gQYssX/v8d8LLc8WkEKKNvwzDLziSgcN
AH3SgDNfVgG05g9JkNlUr58EWUUESVFrj+s0DlBwRTugOlGeX8xymLD/H+MZAOhkIOTVIJqz3DU1
L9hzthK1Mp9I6568pDRsVnw9MPZqZEkCkp64NensouTeRV7kxFa9HWRP5EuYOe4iPiK4LpqY9pZt
YI5MLvA7pMK2hkKQ1ZK8rrjsnZNaiutQ23uuDcQVInBM4wEUe+wjyZm1MUkZFblDsiE1qBL43RAB
b/Rr/vZfVZUaxe89dMgOSoQCTuFTEfxW2QEp1SqyezJgaR8aAo5BghE62I2EIBoCq5nZs0/L8uQI
dL1Nv8FeJwyVHCg0iX9JMmcmnluxSTBp61JTDv9hcx/Xrx5fw9SnuOurRc4RbBqVC/t1baRWtpe4
X9hE3oUsFFCwo6oPotb8EErpY6AZ6QvFJeCcfjLD2bFXU34UrEXSIeLMUNxVvxkfghO5VH6kDb08
L3ofNnyCFcu1scT7NQMnc/TGstvFtfkdZz4ZQNVtWwYwnoUHmsLMwPDTW7B/fD9QKqZHiTHI1EGH
M1rAVe+OQPKByt/0qZatIvl1EyVDHyuSKvXh7O6EaCrhS44IzvaCXl3U0KjrQBTJgaNK5ivSl8Yl
nKnZ4QT2JpzX7e5gootydZu7/H8y4z1AqKqAjXMBaFnzqpBus3PaUOiDx6NjJdlznz9v3TGuZV1L
wllGmNRx9Ae46RLZKI5ayNMTClFT6xAKbPa8clMUWPLDNC+x1mzVyuaHmbDFn+N/XCdWvU1fMdYr
CyYz4/fh+d4G/GDGd4fxauAwLp2mexsRYNw9q2EMC2iWJpy1hRLBKuuXBffrcMyvtzaMuVkGlFVl
IG3GRrtkaLcAO5pF9r9/bSzufzvfEn83y16RjdE3JxlKlHPd7vZTKZQmOtEcyc3hUIcuCeWLlCx3
TiOnJkqzkb4qtemLF6y5U9IrLeH73LoJt7NYvR2jMeYnFWYjA9CJeT09KrRUV2hxpODy/5EKtcTr
Ui0nlC2WuZxhywHqw+p3OO26U+0uIX6ufxugkg21v2YgkL6NFY/5VZeouCmXRteLuZsDwi6mbz4S
le4zFJSz7MgXXnPNY8W12p0DukSa5d+jqKCrUCXTkfQfTsJGH73xZyv9uAED+gx32v5ruzDWAAzp
n3ZkKQbFS0QtS4qI1xQaUchhj85mYUuruncSVOa2YXAav1dO8ZSfoX69aHLvLeBiokEvL8tY7/vV
6yZghiDV9BS8Bw4BGLisPZDKJ8BT9xMEvBmzhwD+lovdY4Q2Hwl/6nXtUFTdaY7W9fmHLagcUQ/g
dMNp4676lNl2Ot/48h21A6Wsv3eT5A+dId/EqueN1Ggh5RPgeZIC2rVOSY6b2r1mYKD97cO2hcs8
sAjotuTCwPexFachaQvXQt9spGOc46w7OkPjAvzNccd1AcoZOSATpXlhA/dACKM/qGJoL6zRReZi
qINb4JptgVu9n5jTNlatt1+w3kBj6t/QsrHxDdKEp+pFa8lrDu5igH0bBEL0zEFw01A2e+5KpQxJ
W93gYtTioOs07N5IgAC4w+zmAkQX8SLro/4VtSoJeAWC8hg34m/NdOXBATVnrqo3hLjTo/w2+hza
cP3Hn7n5ZSEyJsByg1E8kZKaMz5S3ULW9utN8eUpLJp6FrZBfW6uAsrppVY9QTihC2bOGWtL30a4
fB4Nj+7bwM/JC8I05Edo8nlZOZ7LElE5gJREIHkVAptfnHwubJpaY06xi+QQshlKvhgz7gkaq/DO
jVnvUZPaF4aUB+cG4PjzCdR5Leg9CS7THQh0BLse5MN8HjEViG0QSnM/jVFplqI5dM8wmFptYb8f
AALeNvoaz+ec3jaZCKV+8MxwxPh15ykdbaDMtbSVk4nIOtxgaqmDxoEJVFT5sWeNFinRlU4W4DkD
1MQAojrjzB4KBLHnjImNSwakMIzzWx6Sp1m+WEFvn4xB6NpHuu8QfHLFrObfoFPi4On42TNFpa0l
C6Q2GChayQ+2BbUw+xsok18F+lfiuz2zqbK/p8tj0pbidXao6yBCvE8YjnBy8xeRM5cZK02jSbzr
xtKIzkNzdgD8+ms0CAGAnuUt2XUsf1X3OqXvluqose70J+qLvv2LaSs9dwEv39iGtQH7k66/HwYQ
jbl4ZXD5ngr9DuKlmpsbVsFmS7nIPRApcIRzKwoKTUPkllqC8N6roMFRYbghBeA71dBRZJjF7mmK
ExPiEmG2QidRVDjJIFluNDO3UPqW1sC9/Io0FVVwBFKHypVHtKMwJFsq9+95Bc3p2nCFzAC2rkZF
vvbFsoujfjLGgbSTbroSqspPDwdtBaW4sF3s9kCs8jel3+o8nCPGe2TQ3gPObrr28s5I+AH5gLIQ
otE271XySfsl5FR5ue+Of3NpyNtPrUk+Ur0pNWkmmJ9uo4524EkZZTyWToUcxcD427PXSjb9xuEA
xIGtR241x77Sups8g5+6N29myGz6cPunJAbCg5sbE+ZPw5PpvDRnwKpnwlReObzmKk//i+eDZTGH
Fb5aF4BC7XrzQlBoruQk2QD8g+619pFFpS1rsjXzO+nc9xJ8TKO27+U8h5+hB62hIvHc3V55KZQb
5pjCzyAIuaQ05m24aUQ5HTImZHCtaSsR74YkmhZVYuMI7N7mxTln40aVUv197RXjCvI/PYuVfhmX
9s0X6qkGxDaUbP35dlUd+DzHi1+zUQIKr9jb040uSlm9fK2hjWEYgJrkaenckTvmRSPFe+qjzc9z
2zINLSAsALE0xc5dgdoxWH/WVJKM/+OHz1m9FhEmJLWPsav3plhxc2YVnnkz0owWmcZGlx8GZdlo
41DOhROTmbFL5jR39u7nGTb2RT6vCWoXCIzbydkqUAt0MZ1XuFaVZKEjxKy9CS6qaT4KBsr0VH3G
JjvM2HYFMn6MIcyLZj6KOn/tHI6/A6XUSD8HjdOXf856ISTEYLstZSHseAhMtT+dyhSLkQjbtDhP
Eo6qqJIrhHEExIPyqdcp2sNqtmVefLi9Wqvz+VTuJW29EJDROOAQBtO8cFyQXR9LfFMdxDW6xENg
TCSbw00Jy8MzXlTc/kQE4m0kvO+bR6aj9LN5IH5uKzu4qBNvEMH8+YU8ZQRdo82ash+yYzuLRtTa
Bz7FduNYHf3ubgv4Syg8sr9/V0876AtHlT5HqAtE2amkWBZCrR3jnEpuZwX3Pe9iwNwlBSfEx4Vs
WR4KiHjlNXAqGAdySuVLA9pc4/WPXmToV1tYiUeAklulISb95v4drexg2L/ad7e9poIowZnr5Tdk
c6Qeust0T0g2w+c/+VSJOaWMW5PrhX+dlhFvuYBCcbdJ1h788EMQJnTqXM+Eht6tgSi/NFxJwBlT
jKFn3oSqbunBYZMf+TTXWg4PAeuiIVLGpfkzUIVqTJwSpQV6TUnw324GOrvlsmj61eUbrQgUx9mJ
nC6j5tUmvO/p1C8C2wh2Hxll4JoIYpGgUhjjFjbLUpUaexXypDQAsS1boBuKq/vbaH/ewvQVgc2T
OPVV8OnH1UfhVkYGF2I5i1Plu+8mqsWDeyKerF4ndXGxCZUDSRiBJf+pXk2JiLmh9+pdVl4kZ6Do
1FVPr/WZ9S3rGvn3lWVcn0JSQKYSj3tVXUfoQ1GnnDFX20HiYZYnO34pFxMWikQGJvYgmENBUn6/
RD50+iyHQ8aTefv+ncOJ2OqIt1/EpUN2mxK2hqK7hdOPhUzBGgsSFxGCvP7nxswSf+t6xFyGatCt
CcFEU4t6uJpJz2UUGz0sSX1I6S5COo3VSUdBKWy/dtoSrSFDWimWsy1j8hx0m0iJPC+Vlcx4o/6M
BaNVsShDWHuEnxPLjXI87D+shKa6ITUbuqLajiPAMFl/jr+K1XO7w+PZYwYTS5iupoJhdZTuRnq4
+skgUv0HEJJCVQqE8AagdHtY7A4lyYIBY57hAy/TOyib6zhpT06OCaifbtr0hsiNopkyJ+cNfMMJ
FdcFqtchl6K6cv+KeCDTvvYVwRgcepJW7OEq3vyba5SeBhweQerwS4lmQ+s/SGVwPSPddYLosWSQ
wJ6D90iLjI7SNYAw/RYde41mE4GRCxWRrRjOplaYpSdQbicW1g0OCqfJlvp9nUrkcqjaYl/KlvLZ
XxsRQC7kIrbIja9mIlPwtphO3O7tDn6+gjJB2J/qBHDr8Kf781rKJ/pOhO0E3STnvC1gra5DvSJj
xO5Ckjzo/6gphOuYWERLs3j/T87eGMS7tcPGLGFWtPZsUM26pxH7kV64vFK6aoYvtlemoACFe67C
bTaedZZEo/X3ze+beildxIvTKd7VY1M7G2SXEdcez/7H+Jpk+U4w8olxAtiWQclRoKW37xukoIjK
vLBye+LcfOcBQ5C/Eux2ZH3NYY//CID8VHNPiCud9tEPQAEmsiSKlEU0oXlOgopZlSvq01VYbKt8
mBG7Fm0R2JIIPqsi7OM4dK+rDQtWtks9B+aNns5hPZJ1jieQpWFHfeRTiuky9aeFy7WLu9whT0f/
KWlMBJNN3zUyLvAyRyEItOczK/e+okaYKflv4+pdMoiEMtoyLaHSREsZGnuFBACu+GiGCngmJ/sG
RV8wZZQx5nzwaek39s77uNw0T1xl6WS0R6MDo01i1fMrKb8+hKySZAngvRLnxV9nhs7M/rUrBtZ1
jgOsP1WBKRJLhWse8kcEUS1EHoR7mPCRb7vyUkAh7TP9VfhMZnoXjNAzE1P2E54AORPWiZItV71d
oieoRPXVehdSGhhcMiJMneXUli0pjqhb34JbTjRwGFCnUItu3PgjyLKzg6P+AR0SagwK3WK8qv6c
yHdYRQ1fxj2gJfCRyVzwXIhPnezCEVb74dWJdWSAI1FPXCj/tBJQqJizihihL5VubqSs/jn772ap
WlCQeaY1+1xr1Ct+oVduV0AojpU5m3AkN5rSUSrU76PwFrTR6lcK1CO+LB9AUIsvVXoloBpUIgDr
Gb5O4mfsvh+njXO0t54WNpulvUGEdGvDDfdpK5H1j4+ETXxYHZjEJPqexJ9/QSRWAPdjQXR6b/Cg
yUkuU8/2WJbCcvBnNwSLBnq1foTceu+Oykcr/MUdsGGnz04k2430em39w3QkkKFfMqw+Ufc8exki
eZQzlqfo7pgH5dgAfpkPp2jgjWkK4KcjiBHrqkk0ogHCMs+aEKn7Irz40vYD5DS8YfkyIz0gzveV
DtWRLnKSFjFT3WMRlK5qccgTKo8XbbGMcdgkiVU5mn36O2A1YlsBq7eJ2hE4kkDSfqnKuEFi9lvQ
lzP1NSDK4WrrH5uby4tc1evx5e/z83OfGzkBYfK6LSQCYJ/bquJFpV105o6qUGwpZJsYuDgSMZ94
o7x9sJl5SbmT1u5nv3cGUuZkhdOBfafZuOYr3NQW8Sylo73MZAr8eUHtkIvgQbU4nRjhVhqKSJYa
JkDxQCoybSEIwl8BSPNqJ9AEBwrSRc7w3LS1XBtAXrlF4wCVhcgSBiCQCHgxtFrGfmzKf1d6yDiQ
bHzBDn6nbwAwWvLmidllkcaMzQX2JH36IgXgcDGFPve9AKZjt6jWAZ68L+Y9MXdu11Uf2Y99xpqt
CiP4Kr3s9QLNiGGojRTWAuXihJBZBO4sYgorH0Wo1BjwIV4QQ9V21yFXjI0ziYbbOEND+BZoxBe9
cSo2XxV676byXYOLagOohO23NQy1t4/yN3TTIEOeqsr5EEv73Ub1gPTp5d2F4RZtDEvHhOKacIQs
jUUjEpLokC39KFA9cS9A50BT1zuWP9w4LBCgFIA1kvbGLnX1ZvNGfT3lORKZwTcAVGK19vELOLab
a1n6eh9CSwMx9crm2F5e8wUPPrgJdKiz/gOAxP23dOThuNxyEOJ3vog2L8KUb32ZDKGZr8SxJYt8
0FRX9A389lNSve358LYpixMH6lk+yee3o8CGTU2qV+PEBj6royaCDDyATz5YIk4QYkNmZDfcW1L9
FUJxmN7ITL4b/RhwVX+n23Xxvvsb1HfEHM/Cs9j3SlPKB2P/aebdWVFx/1I4TtEGiNbn5JWuy1tO
llp9B7IbOM4hxr0WRpgAU0nyl/VH475IOYhQjyigSMqvpl4Z0Fdy4EYQj3UkKoUj8H5XBGzkt2Of
BNBqyB/KD0Efn2ppQtqcL5tyGXjpHPhvFBzqmaWd0uAtSu5/WuOmEG2TeMXrlaYIsBOmF1HAg9u/
r8P7nmImDlowPWmQValLYgBsd6s0gKjTfKiXpcWBOetkWJsLThOfu7asswty5Hh3JiK05lIhzzMY
Hon9wyHHtI0CnfLsKNZgIPY7sjzyETuGRDoQq0niLCmHa6Kq/dCa852ZFrDx5RoLVD06VB6HSbxX
32UUQKPcP+t5J9uMy+sFkU0gbs8aFDzpUMakWBuARpU2jOmhRry3NjD6nvHVDzoae0dWTyvHEr7u
IJ2mqD+upYicX1kyi4lJ9NMlrfg+4W+0XiawiVOI0w2J/1JOQQpiIPqEExXS87x3zUlULAVFbGvY
HHXHdMe+twMN9x0l7+CmH3/EMQOw4G3bGiOoEUaalZgdNedNw3X4C8IpaALQJlmEItivrr6Ljj1t
aa3mYAEzRGYx10mCA6s+VFC6+4AVqAMjpKfrcwn16D+cOnJEqi/yY1bf42BKopj6o3/WSWQzxQFA
CxjInKiWksVzZ/V3W99JI5JLb6mAdAM14RskylIXQOXwm9octTG5DFSub/KoFbzgRxfnlGqwFgoP
fUMusW4YyHJ8kDZ2ejauKiMULt/kcUzHlOsLJn55DNJUk+uXu9hcGOcOheFLBfGoilnguPM2V62Q
VwHnBXywkUlu3GIsmWb5C/1JtIUG0IJc5o5OjeY7l2GfNvSWd/NuRnlWbIFJpEypSOAjaxL3Y6CO
l9GRWikbkl8OTdfU4851WfNnpodwIriwREE2Blo4UZNxhe7TIjxUm1K5qNo5BShyyHLmJjgtBwry
Sm5QVp0CJ3qpkKLIXq/na21AuFjEJk8YFJdOe6Hqb/BpkFWLCJyN6glujPMsg+ox6GAfPjOdXI+h
UjDbNuPOBgPJlNnrcEef6rx3dG9nICWKt//bEQct/NhPBDHImfoY+BNvJI7IQD7ifW2MGn+m7JX2
CRd7aUhxpgeylJ3J39piu+7cwfluafrXOib5Nvx4CvU/A9GMqgYYNhpbFrAK9aPJeDeJbUUuT35N
xe46C4LU/F200ybqnp75M3ZDWVQ2USa2TSguDhcP2uJewp8fxEKLb56NpXrTUFeAsOxeBZgtkXqh
lz+tgJk0Dol8m6kqlROX/0vUEbXp2DbmRYKesSbY40KGbnxiRnjgyoWxkBg9eBoz73U1TXL4FMf7
3u/Q5TwuUE/a8SUFcr2v6JrPzRx2zjBuSMXr73NtdtM+dND/rlm3GubgvaMlGUxQx461jlRgOJTm
tU30B1tprk1NYz5WVm/qfqrAPSyYpBnuqPUulUO8TKqUkza7YSStsXWAw0L6sp1lyhAKWMsJq6tt
WbMmD991IRxLbLYLjshtPRlfNaMQSWqydH4Y99w2ZOU0Bam5+fWBQZ8dPyRQ9cvSr7Thuo7RItDl
oiTh9+/oWuz0JnKtLYJGYvbY5EQclzHX3DcTRTFfY1J6t2DQfHM1kUGlTlSgRTgBB5ekWItl0Hh1
pw/w59tohWQaAA87sHw36I1wKKuabIeN4cfEz0vl4Eg6lxusQZnzxKySa2FP9fzh0+UBq3fm/y7g
QGoh+McrOvUa+fbXmBSamL8rDXym6WhrhVhWJalzBxwzUxmPvpp/7yaEO/P0JxW+PhXFf+7m1iEd
wZk2KSaVxWEEq9aG44YzVLaLwtfCYsWIjZFxj7ihtbQKNha9vFmWj5i32azSHgvZ2mhd3fo8nff6
zcbGar7O70t+xNpj3tP6glFO/fiz51UlsH4pT+dAG8GEJAKjsXEnaLqKJ0qLDUGNKnZU0CD2wThY
v3oPL4rJKjZbw0jw6/IUyNFC9KYjKv0kJsReGB6o2tNnJXvcG6aU7LRf2g3oc2MDQ/swTDI6Dpb+
l4YBRX9G7A9Lt1T2YOSi1NFOmM6rJWmORcHUUUsqR9iHSIAfi0OEaAYgtr5YvE0eS7vT1Vv3Kqo5
sWZ2ETp8Lar18vT715xFA6AsypV57GRJT9RF6b5N2k5ezE2Z/N2HJn2IwVVvGTRgy+EJulYrRUDO
tGYoo5xr62uMW4+9YA/M9Ygi5AinpfhmCGZi39r562ZTGMeeGDCQZ58hVpoISNIZD7o9UYKEkf3A
zZG/X+bwxKdGxaCRXHBM+Fa+GdIhskDNM1joExLaUMTvlVaxNavH50uTJuazg8LeOEq2L6cseTyg
Jk9fQlzdnQOYXAtQdejZCrcagx/+NFI9JMFv6GK4pYCHCqkZUyopiHFNmRwNq+GHd3tDHzLnTYV5
OTheO8XC0FJIK3R2t71MpjWUejP9ajXJYjYkfVHHa8CAD8VYA3rubCtjhSV3u34DCanpUAUR8wb/
oFDrDUwoIK3UTcOLWJFW7ASqJs44PS3NxGlRy6qgJob77pZKbBMs3X8Pv7HB+PeqhVJ9WFqBdmMD
Vm082Zf9N5I7BUCk5shOYGGoqAlqQYIbd81UJHHdENrXhcB+SLaBTkb7TgfzO19/6SKco2jABtv5
2SL0jcKKqxaaC2nk9HKDmOcInovfHV4F+tRbYPbyB/5okc72SPce7tCewhQ84JE9S5HpFA6036wk
SZp0ZCyMBzUZSzmFdMd98EZjYu+LgYZFBLo/a8fsnZFs+B5vUc5znUnxefuWUF6d5qKHeXKqDBsT
KLWUuZsNlBrIROdJA1lxE6ioGj0nc5yev2ejQZ3GuDNEH4aQ4yFOUV31ikIl9wf/p4X4qJ5kk/Dy
Z0B8nrPj8mTF3rZFhTlFinIcKZAvUStD8FUNzTx8VgMKOJy9qB0+Unroebrhe1OkOrtSPIiSl297
LR9ExI2Pig8IlZj6xl64TZ7toMXMKVYcg9r0sKcJbktsVDEMvjwKOpcQCmutP51ug9uTa/T4txO4
OFulRpIlZNqMPWW/CZpKo245EOKNsMOH1KGZ3yCWxHYojdf0UKneUju4mCsROyUE9yH3H8OStlgt
Kojh7NmdXrmAU5MshG7sYy0N7Y8sH0FD75LvwDn8eeTgmFyYpoD+GehPXLXozcw0IgP6t2zXu9hb
5cR9PECuTOuz4Z+BHSBysoa33lTDBFUzDlR79NsBD3ca5zS70xfihAoy4i0no9o7HYj9fBh2/JM4
rcnENa1Mrrv2GAiZR/Q08KYpmKAJ7WF6QCp3VeOzFgPOG5wku8/HwdkOMopxZpsT2S5Lco+e06dy
OIGJBCM7bKMU0y9X5BLBjLcQMBbWv8dlJL3ds01rHANzS/Q4jSECrSTzzYRKO7NVC/lzZQckR2pF
3y1tCew7o/A2qPEpF+jgkPCnuuDuYbiWqnPAnlMF4kuI7cNaezMTiuDxCkY3vclTAwC98V2yAHYK
HE4mgkjl6XSOXJQDfw+1z6cRXLwQ4eHmqARK/KA+EXKWxV08CzuPXXvaCUtjLRyOA+U67woftlYr
t1lk7gIRaF1s53hUpy0wqHKHyQn3L8DKXedeiQDoknyV3VhZ9/zvayvvxiQCC0iiT0bRGc9rP98f
SzVWsCDc4X5p2hmtDzNqaRKZwucxNhReBCkQX+TrybhlYZwdioKP6Ujd1tm+VkZSvurzzumY9KfG
gzh6AQYtDVKrqGraGGs5lC5+LjMEsF0UsZvwd8+04/276ghoxkOlLbpYsl16T5dpZdufx/aSXmVS
h6M/MTm8hrCjEboA15I7z1bh9OhJqVFtUpDP9GQJekbdd9+R14iYT45SWF3Qp9pxh9uDvT8QNVXE
//OJhGJgmC8Vln+DVljqJ56DSW1alJQx1M7NcGwB/g16RgZlGIj3VeMoyuWib1Lz9TwbV+zfeLHY
qJWIjQxknolQsq7B9gjXLOa/WgxvEwcy0ASTDlqOn2ubyR9tEZlDwgAPNSUzN+olEN+DGMijeZMV
zuApNtq/nq2Jdqh0DbzZ5liDk9iHRtS+2Y96atlYeqFhBcJCIj7Dhr98GDHnn7MXWLoIM58Ilujo
bMpLUanB0pfRl8h5EqsBSrr4edhP5qpXZMXi5rFiocMMkseNuSuwVTIK1dSFCAuBGol7wbDBYBmg
QqOrv84CA7jJjL7A2BqWPb/wP9RW5N0O2BpfmQ9cvCEGifqPNJrN/gzePbwN+NSzlhO8EywnKtN7
pk3saXjxOM+mbxLnFyg9x3+tzsusXB2wI+fqUFWcRdIoo9/E/aliqAZMdHA7uW961TYlkaTLTqt2
7wqh2CtXGOr7sKiQIcr+o72ie4Dti9G5eSt/nOH85kquQCKIdTKwx+OCQFjaQN3pkqqLNi9iLnn3
VHyITu4yTFMew5oLQr+OL7C+49xsYRxn7mG1RKRQ5XiVki+1KN9Pl21sg1KryvQITj9UyDpfldUc
KJunyt2gv8N/0SfBUM0QaqnJ/Tmpe1w0hvZuiHRaL6aBIZxRFwCAO0bKybgBTAZejr8clJu9+IbA
yb2SetzsVDsL8XkXzsisMIqMbx2PPjaZSDyqcAC80vaGaRUQ9jwAgKK5dP41VKZ8F5Iws/IBXAmL
MTlyVUqzYHA4d+mLr5gRp/NYH7wRsZmGPjFbnI+Y/elcHxW2Mmojy6oSk3ikFtc8ak9NEHBsxbtE
T8CQgFVqHAQp7hNMsC+zF/1w3tjSE9yByV00vdcUmbxLRYy7RizWala3LABlqx5Ejj71y6IAx2k8
WL6TQRRUztLksgvrn68jkieYEpi22/mwmcyBPUeIGrpH57E0dVms+YgDcGofRTuD4zdRLH1HniW8
cwOzxgt/dOftwjy4Jr2+4fzJYptlb7OVCAyHNTlFnN+aSUKO9EwneMk6oOg+nnK9phrkbXSubmaG
jGRH+1U/i8OCI3YCjjoZx1B/kqtK0W/omBE3a5Nsx7IlPzGJKTheJSZ8jOfdtxlGAbwD/nklwUKU
Ay22eG4phhu76ED+mwZ0AD5bJ4Id9gXAyR6dcccn6xkJTKeqRut8Iohs4UlGgqQLwDW8icI0UPjJ
ZU7KCVzoCqHFXh3KLGVdwitTaIZKFtAy4oYMUZ7IgwoUeBJC03H6jE7mndodWeGwVcS2WU06alt7
uGW1wC7xRPRCf0AsT83XVXFeOUMF2AeQQeR9Sl7U8L3ROeYXjfnevIWy7W84GHVbg8EBoyrGoBPQ
XwtJfkZF6W0JqfC35YuhF40cbS+L+ztlMijLP1q/t9pgrxQ1lgiahnLQNSzIn2SI4afygL41GN8m
I9ptahNpcfR1z6Ru7puuiWqK9tJNnl8oYpW7VPozih04qdGeJS/Gfix90ke/t9vfeB778+WwZM0A
ct/vFSilF83Ht3Df0mmfGu6fzMuZmInySbpZ8gxQ0rFZL0rhSOJOEzKBdIbYJHoqHJ7LR0PJCs3L
e9GhAH/msCQB70wt92fr53r/78f0mOS/Ci5nz6wUlmx7fc/L208YqFNzrCODMVfTky5OezOHcyS8
Fa52R7bP3Tu/EmJJwjMa0q0MepxKuAT4okb0eyeVy6NZoXc3vN3tKcbu6tCqbVzVNQK81TdnbB7Q
Lcd+/4aGI2guH9aQWCru/t9VOuww4sIy7Ysm1+FOWGZesaqWlciK1Y3IWpz/CB+y6ua/Qc3j8ojE
fKAnG2zLfAzd0WPGNukNZdWK9i/yhR4bEsJYr5tQVlzgYySTqb2DsgQTQ0vJYVPV/prFO7uUFuAY
wz/RzvioPPOdBuYOgV4udmNtRXnpAfCCwkkfLdXyG68l+fycAW9gAFDRfYSa9eu6FJ1zWpzxdasr
UawV5xKlE2w5onRNik98dGBDz/1CrN2Ytpob5DlOizTL3WhIvHCA6AB6eJdst49VSRx2ZwWt2Vx6
6CdGHoDYc0pUZNFL5PaO6oyj2JpZRKfxrDIK6dc6FVOUqnKdAFl0gmztBNyQ1mKry4IdgRYJmmad
F7h+plml3jiOfDuzKDkkqdiWVEKFugHgqp+uzWnpbEzYGnK2W4Y4jfP7Ppw9oFQELU7LGuQJ/R/m
GqiMehRq4H5IbtKiL2aUgFdRKFlVfEnkIbR6uMDjocJogTM9UIZxXuM1H5+edv8dcVLiXA0Qw3TQ
G9vinZRmnyQhYM0creyKxSSLp4oO03l9Jo3gHBtbbvQ4v731jPTZPQdAhA79hAplUN8DsaspPAH5
1+Q7atNvyTvKK+tlO2oMKZ6VNVOAxI518w9LTVayAd2v7CvLhZN/qORKuhbapNqMSK4xdBEESv5o
wdIllxNtIZmHQy8hKOTB4Uc0cO79O4gTaFGbR7fztJEpAxAWfHND/97JJhW5FntJ8q0cK4JgDBGi
WLCObAdR2bOsMQW3xUIIDRM4TVlkoiGXPtC4MRjpw2e2rKdGeId3G+2Z43KJnslErBPPtsN6xQjO
cLU2z8x7z5nn+SgeVaHX9FbDszFqahvHnCRBz/kfLXCiB91R+4lKPivIu3ZzdVNunfn6VpK9pdej
4/nQADqXfPZ1eo/4z216hH5q3pokW5XnDMidXS4iS2ULcVPRFhOoAdgG+TxnEYN/xbHIrci51b5x
wdz00R/RHCzsBDWEC15hcFVW1LhI7+cJpMySgUn678I2J4KsnYWPPfSTTtGGoLxefF58Unpf+RYV
ufVArZBmNMefMaJU7vr8nNjdsnf8uYXsc5SR2jWvBsMdzGdrLY+kSP8DzrKR754/UcNYHFTjVDl8
VmK71Ca0ETMErUCdxaoEsIk9xkgEWXz/z2tuRWoDj0azQbC30LThM8/3FQKeFDnaMXvafZi8zRHJ
6kKzeTuXEYOU7hMcjnq5VA7SGoZtWHZPCi6Kcv6eQvWtD4mYUZxY3ujdIgIytOllkmI7gQdGCOSm
qG2PRphDeHiZsNdwLCvd1utodN8rsGUesbruzFS7xSQP2eHdVSwJDatbEKfCSVOwaCd85l9zrSQq
OuOSLhexe7GqRmtLypeBVpFonrLLY6PGa7Ip4xierokcPNJ20JLh0P1yF3os6XwLXMdUS95Gq8yX
dThiGjjnpLjyRmtRZYg5wZDXjdNNtQSmzRgnMSBjMg+DpVzcyngHTgN/VaxR6eREp41EQvJrQ8AY
MxqMKKSdr08OQ72kjdox/6zp7vH/LLvVQPnG/3E3qLuF+aygoeKt/uo/vd/ddNeIuDmmMbR4TfSn
E9+OlwgMncFfBf/2cS+Tz5VdX25nhTHr//0/ksI6CQKXogtTPyJhx/FD8dg32rcsyAG6Ioo9vi8O
g6L70Dx4V4rV7ZAOXvemXaFb+0szEx7gHVpV8JvFmHpRaNjuxhyo/3ix6trYIHWZn8T/KdtlRJz7
PY0yIM1Ba9Ip1Ps5TkP8WPI5XJ65vLRTVuY6KYPwGrN7R0/ALO0oipD0Z2+r8D9R5u9woWzdWISz
AD/iJ6YiZ0fEcqx6r0edRkDLbnRK1Prh9OOf+ainis0lAfdWPNN1j4nAWPm3vBrfDr32lwXjpsVs
k1pofnL2zLV1AhnfOQez+0ZGjjTzDCk85MdlGd5jYqZqa4dAd+41KuK7XnISpZPVJ97OX8nZZhBi
/dSeqDCyXD0wMdii14GDwlFvXj1d/v0v2ThbYHIqqhEZO86vn6gghK3+k67d87vNih6z5ASS/pZd
+ItrLbBwgXypr6qOlGTIo/71Pj069CkGF1s+1G9rcXe2oKAlrfN9fqKbbqMidKXmSLkxoBH4XYrm
ePE/dMsy9mB2x/h+m61o9OaINpQvzZkBqhFN+8ipt6TeJKdHdxQvIIsSrYIQVG9ZDf52E0ICooYM
Ed4DCR1jXciCmrkfT4zXH6m/4Mbo0vCYCvUP/eOAJaS/h8J5/DcIJ+j08x8+2OgJvmBTe6rRQ1oq
kKLgnGVt1ipJFR07PIDmvutEJVuwDrhQunKeYEcmLDl010G39a1Op0ImZJDp9KzYNMe7m0PAtGto
T2MA7HMljnoiQG2c/8gpeVn8/bGcJxpWx3zLSF4o4D/KumKpMQi0NLiOFGkqJ9wtP8iA1jnLlZub
1ROjTHtPN2hfbKid5aZ+iViM1EeIADmVN6IdiaRF/BvwJ2ncZTb38+LNIwxS9F+EDHvyvFm41N1/
ce/xxoYvW19QbN/aox3p+rtzI9zmBSW7oLfc6X45PbEYJRDvd1EBVIuE9Dwglt6kwf3M2sY+sUmI
kQwF/U6i+ktB6h9UbOsfVf1M4dimUGNb82Ff14T4ijimuMSjpcKzlp5BMp+nmTsa0ph8PGOOV/iq
titET9g7EfmYeRSh0F/i1o52HJ1zmW30sbv0fNIPKGTukZOoWAFD2c8UpvW24dKYoyqOAGPQr+5J
Gc8ctCYS8pLJwor5vcdI9HEyA+DRRhvWWG1XqGDRP00Ms0Q/xboKTu9OsMwjLibF41Lag4JPcgsj
fCxBLWQeVT0s+ZDG95SZ/6Jll6XzoWQP2hkXAWqicepRGhWr0dIt9XJCF0WRSWn9Qy74S7CevWrh
Kif+g5sLeXzRvXO5VTOhH+DSYVZRionw1x/jRvObfm4FJJyNqkIkphZJNBe8DPTs0f7DMOaQhu+N
bh35ZCDAp8/qy/VkK0ZP/92UOiJYHmvNAe2ONnkPRM6ZXPhExs3eCtJp+Qu2bMf+OMrwwC66j+Iz
gGDaN12KJQEQovCy+rxgKWautB9K+ta13zKItQmbyUw7bXWEg5LXsb0UKm4P44NtKzEdjQyzY/lS
+jSuJUp8gL2oy2puL5cjjrXIKqPSnYvRhNpsCJYgJwUJ51h3Ks5YG9kYU7nWr8p+9ovlzi3soNzR
YnlTVQykSFZ66valdECiAKtGsSockwaIbnJR2x05PX6QYWggVWNWg8RBqEs1xOd9paEUULKOGsno
pTz84/TQDnwEn/9VIz8bJ98Eq46IeeyVrd4AuTPZtma+xH1VHfmwMQR3+EaoJDZHeP3PeWP70aDi
O01JwLPLG+ORl9bpr3719pa/t9HFIysxuzWpq2DOOAun7hn6hFVtr5A0U9oR/nDBNWibMXJNd8h7
4P5KCdMc0G6eAOZDA7x/vmhHocUdqEgj2s9Jsywn3/A+jsldiZHVp9ig1/n9Vyn5lxpcWszN8B1k
OOEFax/BYPkoZ/AYOvn9i1eXWFLku9zJ4zpqQjDOxKyQF7xDfKWW08bxegUyhGms6LOGTOCJxhzf
jKc58eaBrrLzXugLKOyLXuKIDoP8Vg1KSvh45aRZ9FNdsSj0TrOmfKMxyLmbdtD+LLhiB3nkD7uX
q/CWcQlRW+CMufOmxRJ4SEUDxzc86mIW3Iih31YwPf78FrOjwLET3FlPPUoJAVXW8RFlZJAZ/ytl
FYqYBrChcwRApzZfI+rNhBN3fdXZLYQU1gsjscrIcvS+dQpi95uWYVMEl4+BdwlhBc1sBSAPHnX7
7Furw+0M6jjIvAMli1nGfQRlei4ZvBEH0rjWewaH7DAWgAzWuoPsPH7s6CL6Im5fGJ49W2fXXIhf
ogZa+R3RhS01+irwgnJcX06t424P2tkJHCx8mMrXHkUJzqLleM/120SCy8GF94/lXDSfS+BWGJz/
o6sPUCzGpMgJa7LIYei4ywdTo2V7N7fvRCAy33NhxCEk54SIeC//cB3vBqaG9K4ml8E0UzS8VF5q
cJKZQDEdjX3Bs0bsp+DMfrauLNxXjp8z/CSx7n0tkluICx/TSyUv9QuoXq+09rCia7tA1N050ZOB
LEFt85bZ97AVuDrlhXUd1jlD5VA7n9RftrKYrtWP6etx8BFmZdcUBGFFSOzi1ulwwniLuMgxoEq4
eG6em9SrPLciDXAEqhYFmnhJ/elyvVJfCzuWNU4s7MXLLpcPiOpkhwy8IKouh9yip8vDR/sPVwqu
rgRHBWGQa1xFvXXLY6VsArEFM2X4b71lDENdtvNT4pa8bfcD1plMM3yJAYPvYDfnT4t3R2P8/6lQ
S+mO9wSDCkbEnrc2Pz/4UpJEnTaYnDipAjHzToDsCsv8UwBjdGJu5jr0Y1frHqpdr8i9O+y9b4J9
7oQrh3V22Atzb4kg5XQY6zZntEJgvBRQykuK7F8nadwKMO53j67iyFr3ZMMRh24eVT6Cv4do8yBS
wlAowtVpMm4PSkozn28qCVjmX87bMOMDB8wxJDc3LVPhnTQf3VX5xMK0Xklsq1SNn27vbVcvsQGF
R3BQ8vev0A1Lp323ncVFyzTiZ9WhVL3PKO6g9ltAZdSsaDw/at8Ld9/O11Ld9UAiUcV8EfSEAkSE
Vj/myzAerl37KK4ewkGZO2N9bgqZTO9JVMNHLOAhuBWFSa+97U9YFeQgl1mmKqm2uGNkF4DH62Fb
nOwJ93IuQA5bKZQI4Z9hubw6xkDflI0LPi+mj1gQKWB5pUsaejuszf8UA6Ybe9NoAUm9tqeqgGJ4
E9WQ5LFB2XwRusgHqPNzRuToUIrGkvrpMUr/V9hfjC6uDDo05LfUfJ49LNEN0YOhAeyWSFmtJKCz
YpfiBHQJ9C3F4ic0wJfhJvQCTZcOS9tLZ83Bf1ToCaEJUrhGaiJd2s/qH/Gh0VvACOcuxbqtPZvI
RSup7Cb87SJCBWUbs1ouZeYmIdTgaUenXH6vlDAEBoH6T9VXJ7Av1yENUkXKDEg+UnIZOVOM1i0A
0uA/zTZfSQYq/VxkbTuxEvdKis0DYG3gDIB9h4fgIMYU0vXeRU13EXx5oML24UVs1W3syenZzxJY
Pxbf0DjWr2Wg0CwXhbgmT25C5/XlpmUDeLdb0I/WldwYW/rL1tIEX0Ns9F1+Z5waeJaEDIWUAFVt
QCvW5sICs4YnhfbQQW9o02+5uazurSI4m4jnJsoAgUbTKZp82Z/204Gulms1ibLAn3RGkHIDhVGM
QyKisUlZMpFApQJWXQVa5q3kqauLJBlJ/Ju1WsjspNf7PwYQXwMZWjtnRPaFPupqdx+ZypALOBG2
sRZVRWM1DzM7Ta9i8rXZnaZIsUUX1ayVD4WzahpWfd/FV4MClyJw7xKM+b3E1kY24uWxQv15H7M/
8bTqlwt4s9s69qXbm4CRLmxA5ubxx7OVJQrNXSiWSH9S7t32NAJ5gCZ/EDAoomfZC8CBlLqHbtXS
a7Or/6ZEDOFL76iylwt4pFpJS+QK6iDHaNHcCKL1Po+y9Xaa4Rw3y/rZiA8lyEIr9k1r+LwjslrF
Awb4dEv/BwrFEUjGfB+o95g6O/laQsxlwSB/8L1O5Qp8oFwZlLkhcVycDu9HsmHFenYMBkYxRXsK
Tg2QYtPKuT4s5iRxlA2aJR7zPHz6fcukbC3gV40RD9ULUEIGHo9Y4RaaTd7JSB/Va01OD6LD5o70
nUwmJnCmv+9kpVPZgHu3NKy953wPHi3XMSCGV8xw2E1L08EFxoYgFsWfyx68ATee/7uYG+2z6YxX
tR3Z9nu0NVgyzvu2p+3XGnZcLpn/BCZCxFDTnBtwAJtBMCOieBgeRLjO9KaqzoPF7/O2R7GId899
PoX2ppT1eizCd1TmZaIMFSrjyg+TGqL+KhZy4OwjPQHCNtZO9hzP/9s8G7Rb/Veo9mFpkflhGAFw
oFRKGi3mcZkz3M0SixTvtweyOI3DHp9tdyZ6IvI9gXrfsfhpEEBPWHAmt1nYhK4WScZZUMLiJK8P
2iNsR5Ay5skz7RmHq+fqrldCqXKCUSvpnSKwgyhR3S30CxCjyERY8njakNYqeQrQqYZ0dzoDUh++
Pfm3bbKfDcMIotxfjDb6jzq/T40D+kPWCg0RCpgtjI6/jgX3ltlwz8WwmqrA++bSYbtvkkVEDXkU
qYYL8V/Hp0vAum2AUpujHp+h4BEVt2LHW6XzQ2m2/Tghvijy2lsDHyn7dlDsJmqM7mxOXJOJAhS6
r/QxjbpgjQzlVfcU3DSWPLkyOLRlxJm8aKACVAxZUROmypGmvTnzXyRVlASzJtzn9y7nCeg32w9N
DuazNCuvIO3SZUP2x+BXkm+fDNPBM7y65s4/yVA/ji9M5tTyV10Sd4EOk8ETroAMCpKjQ1NijLAR
V8QW+EOeuSKfHB+o2z1FbJaa/nLaoH7RicNYwPcfKNnjTHYqMFGSeU813/GhF1S4Qb+HKZb+lCad
7SgZT34/YA/7l1dMzt7NVJxVlPFHXGkYr0rtulfgZMbYIk/lcIWHj1uZFMUWa1zl+C7ZiFhaPYLr
0OmU89UNnuvplWoochAbk1p8wZFFn4FgB7w0NuIjEKLOuWvekt31cnnGS+4Gv3e16ZUGK3RQX4/B
2I7XfTs67zzGPlU6yWBZAtOdQEPfLeBDdqTsRYSGcLsZtnBoG0gBcVuCuOHNP660KzbefCskJtXG
IMYkyykoj36OO3yJrpBakrmylr7u8umNvrSewY3FtmaWzYJLmqL9bIVi8mDZ9dBs0+0YI7mnsr28
WHQ2b60XRQsxAjU02CT5SPdUi+NjZDlvxdnCCL/jiXIa4zVm6EMWu3vTLYosPv2dK5siO/zekkd6
9rFCSSB+u2Lb9phetn7GpPjZUJEwXlYFG5NGV0n8PXeAIZqK4AHO5f2F5p9lVGQptPT4OqQhuo7V
i+qnE32RwgzGKoMk5/1BcaMPr0fWPRQ9zv9gnk/kja3s9/giLO1ULaZLDCb9KUVRshXQ/nANXFCG
JhhD+X34EErd9AipN3C0/Mqp77creG5g34RMrjLGCCw4KYp5pXOn8V0JExJxi2TxNMYSJVCrU0jk
YLDrOiwBZvNqwV9JmcvgR38Jvq3yizFjPLiHZ74DPEmxaLUCtky1dEG3WiWn5tj4I6h3TDfjPsTV
pviIJ2Piud6rf3skw9EXNKqxgKEamV+sJ8CnkcoL4RLFRN/kjRQwTuzvqMBZyt+LPtI9bMPu5BLg
/mp0vWYjJWGwHTkhawLLyVeVOTLF1ffjOUt27mByIsXN8wkuaEGYjrTwmWMH29UKLkt+ybHJ1n6Y
2JUgDBjyDPILjDYnjFW86xC3uofzXG8BsMCmCO+mHmsRJzC10I+3WnO6CyQeHkL595TYsuZZ2/HC
XEbeAX1/DfzNuKFcDIyvMAyJ41u4yGqucKhJGLQ5+PNWyk3pz3gYCFR/KHJonQfy5bo8yH6/n+1+
MjBdSudQxIrIw9xtTtoKX2dj1ORg4Yv6iPqt9o8P9CaUh7GxncLXDMxFfQsNcZ2QqDFnk/tHzDJI
2LQ2rlg8FERfeTtYqqKNG6BgFwqHK3/xzyWbh+Jdo+WmuHsvQppNRbdU+5CRAnY8Qe9Pn6eXVrZS
p3SYkb/Wf/NlG8IP9erPsFXpaINFfUX8XnETwHG1/gqr2t3FwYwCp3Ni/+kQVAxdz9BIm6gZB6Do
UzOdFl/CWlqN7xFVOqXYNW1oZRLnVoArci0JGdLjnUuJBTP7xd2g5C3P74oRYYL9LaCI8HZ6QALM
FHBbzgtIG0zG2VHS0+21pu/o96+9nVs3ZLG0qbMUit7Jdl0+ZsXdSCYAmWvh6sX7gagaZLwXH9Vx
QInKPyQ3ndbA683FszhTe6meFHKvmsnYjqWRzIu5v6Yz9Zpk3XvZ+SM1kpTtP90GkcnWX7Mkn9tP
/HQd3b4JkX2Xr9B2o2/RuIgoUOVBuOukRMVHfD65lryOpScfSznfA36+PSfyWR6P3Sy5Zctfol1J
83aKuL0QB4LHmGEgPa8Zx2h0qp4inw1qJr/w1IQlR7paPrcu3tfAF8Hub0O8e0MPJeqVYz1ExsKl
yWArOOUty7XptmaYwidUM+q1+FZVWA+pf9+/ZPxRqkxZm+eoEwiTBi3mKC9S9xDtWRntXfFU3j8n
/AoG9LPqO3Hl9xE+w3TnTsbvUiahOo9BdnC24G1xikajWESuRd/5o1z4J4h/ObBTyF9EDa0pyoD6
7Hacl6iDk8C+3tVy/XwB5Xwk7/Uc5dcfgiE0dDnHDAW+NWfu/bXjIPkfcWsVHUCkDh94AXcjyC5Y
x0M7qOL7kjS+MmOjZDWl0fXaprDJiskxyfq9jqB3xqZhNODEmOPpsE8gPecztVUGbPD2+MhAoNFa
/6S43QacAOcGFm2vYe8WFBBMwUmzTu16VQMjYQ4r5qXoqMpd6ZNDNOz1AO3b1+tICFj7HbiHl4Pc
KohuR9aW/FnFL3ESjm8MuCQRCO7xYrV1R3HAg5ImSp2NUpTykq2JxYY7f+9AXULEfe2NTgNkehO1
uD5W94dEeU8jpMsZd2EvNWvchZroglmk8SygQfim/Dm7VMXSgVROVgMhqD0UsoHOGhETHOkBmaNb
BIK+/tZq4+8thVGZZPlymmMPPqatwOK7Sguf2lQEGs4XNF29ab2vE57APvTy4Ed8+gaH6MarsOS8
9k4t71R7cNUU6Ubb0BaKbNfNp5vAFgsgmh2RuS9EObmHebBdZ2ejmdiQyIRtDIKxEzb5QWav0Aqw
sMg058rnq42bF03WQhXB5zQ8m65hwsptBYIdCTGok1eTSKq54E/CwZCFqDACAnCVGGFfGvLy3FwJ
C2BFFMqmlynz4GjYH/Uc0jtIxBUtPUkGsPRLqK7oU7s9o7g3ApadUnWTPb8mj7ThEkrD0gHOpRyN
tkYA/9eL0/Xsjyg6FChS+5LCEIO9NRJbhOaUCVQyQkY5uKhgBfar8MWizSycs9/r3C4AJPvWblCO
Y2gtW0hmRr7Yty5kkSxp0nAsYur9t+7NBs7os8FYu9OByz/pjek5hmugJhHCaWvZfdU3j2mjQTQG
oXkfutXA+6aZMjZaQ2yjBj4upe1XeKzmzzwSK96V2XzzkXH5Hghs4cnMBF9aKbpmSmqmznqWGvm1
IXdGZXsUGY95FZ+Vh9rGhZNfHfTtKl4GYE/gAA2i4wJW2qUvoDJBlDmtc8HJFjlDeFSQ0bxkAbcN
DTBwimPjOY8h0j9CZzdgW6lnrFHK1KX+eDgiRWMuhvWyMvpcE99L3amywIl6ig8vncnYfBlDxWWV
cKZRiTH26OG92B7PDZ0y3P9Jd8G6tLYKFJJOJxpoe8/PXuymnBXDL2uipFTcOTrQNAhamFqp3GaR
frsirswBIZx6OuocMaAFFghRWmGKYYQne/eKGG2fsLXYaQQxhBf6G7vuWX7oDuBi9BZWC8AtVP9m
w29qVulGkYnDpJBvkirsN6MoCKtOZwYgtCZbm9u0h520FgeIUXEm4NhSSWH6r+BQk/qazVq5lvHn
OhTfLPFlknCMaAcweuY6dszr8i7UTuBBuePt8/4d4wspW4IjZgCEb31WdwZVVJqbLi9Atq9CevZd
C4Mfz2DQVOMaI15v2auZjcQ9+Wjj10KutoinDP9Vd7BfWI81Ny4l5jK3RzlneVW2mEiw2nALJZUp
WuDTT0viDB60AV9MOUUzgd9m66uzT1KEfYEAO4qh6I9dwULxYrRFqWKn3NfDgzO7BMcbdVF7IOU1
Rg2Rp1O4I0oHBsqdsLcD3OVKuFNtwUl/RoKp31e3+2Lg9C0IVoZR87e6Z9S+CLrND6fSMRVzH9y4
9f06EkIcBQEaQHRldXZHHj25RadHLpwGJ2ISCwviKI+89L1lKytPp1pqwu1mowWbyWvNb4PkLyXD
dnCv+zgVssoZXRUP8wIEqeIUYlX0i8OOISzh+1drUoNmxd3PYTmdRrfhoYv2yk9aay7j1lmaqFPQ
llY/27UgKLk7HVod77z1i0i+DsZrss/6hG9O3MIM/zO9C0QPu1vMBIrPTpvzcqIktnIM8/e+Qxdk
UyZzXdJtpiukEyjtAJ7160mPLJB7Mpc7g8Dg2uLFHoODu5HhOm0KQTvJy/EpqQMrzR+YklrwSZU9
0VXtUIvOGX4ys1SJszy2r7y84jOD19bYVcqXchqEhY0jsrcoiQ+gdg0r2PCj5FIzhpxDay/3kPKe
b4Ygi+BGm3WuWkl98VtdVGqpNkdXYe1OJR7xDbaWtcQbwEvEy6SeqR8VpK/W59hzM7UDV2HvgVJ8
wmDQ7ad/1SudG53AsEowtRp1LeglHaz8njpwMjyvNkFTVBGlIqMg286JXGw1n5UvQLOcHmGFUuP/
AlGqxnZv3YqIZIeekgP7mMpv7jTr6FuqSXFD+pynTRm3x0wB3447dnUfCSWuHJpg1Hl58ukHT1rb
vlXSr9umITpFpOZpWnpd12vj3nM79lNcGqMjuNzBef+lnm/Yk4ZKOKfnhBpmXfgtGgGCv4nXoJ3u
odhoFad5Iy80w7+dvmAAm5eCmEEQi0eqqjw013k3yccJdVr22LKjRAUAGlSPj+tz6GLEeNKR2tEb
BIRW7RQoV7OxI7jwJMFVsHiV6PoZJctLWMj8ZgCmqJndE2dy+WAqQ7iRp9cH2GBIwEmSDZpqURAJ
rbwkgJuipPxZY2HuqTZfHVjVPdUvV9t+LnQ5ylJUM/WyqN2QiL01HCU4HWIyH3fupwE1a8BEwMxo
9pwg/v82hzoXhwEp5zVx9eBtQ7gqwBQtYHB2/aXDZeMclyo3DNZLJLlpPSaFVW/3ZsZrqNXrlF/9
TiYNISe+hiDIOwjPKujtdK3e4RH30BpjcJL7xTcZlaBZawsuDPqVTum9svH+9vk3GDhUEXn8Bg2Y
AZn0gMVpMxYOGKg2haf5MUO5uYhSsKjoS06LsLWdEBRnqp1C/gaODo5paFBgTETkKb7aS3NWRxoV
89a22JL5fD/U84e2rNS6QNnSSFOlIsowrbYxxXNl3OasDQ2RS18SZscpMFCJbiZonIzQ5jlbAUBB
oA9CZsvRZPt3JPoRWgCGZ8ma8Cdvh6kKdj4rbP8gXdRqz3nt3H401TbjRHRjWwGj25PLLDOPSHyu
sjGfiMtIvK0fEuY3oqyS9wt5dQV0wscDGpxOekj1CUKabtVmEqmkKAhen1Pkr7NCbGZIv6eRE2dd
pf8aotVnmrlpsAKAeqNS8ZjgKy1BB8vzVMaIMDza23omrLEK6ZlXqhtk5xHhyj3/sn1z3gsoEVfs
XqWHavt49fsGI8p2C/HoEpzXFV6/y7zYM8shQ7UcuSIsJaJCcBzKIYe55AYnxZUs8wpiNmqZsH6i
zza9HdY0Wnk/eFK9G/w/tkWdzkbMNrQwHeTKDsQj070ETJh/Yu4YtGqr6UlSnQZK8ZTY2i4H6Bzr
o3JaWK33o/IVVjck/rr4ZlRezdG23zL3kYX03q59YCaTqdWmEjsaN9ahl6r333H5Dud7tlfP7Asv
xGQb0soRTtWiEEbtR1BFdt8c44GVaWXUJMyWzTdzD2EZndXK/hX8TVZHPX1YeMhb0eld0QTd0iXO
BpbahqEQP6ZXgiDD/AKRPoMWWEnaITAojA12op/7AuwYLUDoI3DYCqfPbUAhQqpAkTuE33OcqduK
sET1LE82hBXL0nBKdagB4g+Qe6TGxuXrOTBB7hHBkzrTqThCjcN5qJMqn8H3kfkvJy6p8tJh7OZH
JbyS2KVRJSnf360v37sokQQB5wVqvbD/YmyWuwlQ1s2UaafbYKm7jdusFO4bmyJ1iBxkOHrMhblE
qDgdGathGNCDHEEICiABgQ+9/IAnWGYnRHrko1Uqz2y7kWycmVUyfuLvrMmOOANFUedww8AreC23
papzwhca9picSFs6/ud8mN5+5C6m+fGJ49pVHu0wtwI2OWzH/BVO5l/yRELCZ8pMBwqNB1Qsextx
Cn5SbzPIApNMTsh9egD8AFiaSTL9bVttBoJ4o539qWGerzhHsjUj2tiILEvd8PW0ZavEGPZuTpdr
CPxinYQ3UjioQStPc04d5fH7tcMWsy4O0e72PerE1wIZ/LL5e5nX/cqv2se2dkHAOWsrg1quftXN
GFlCTymasWNzMRGOQ8FhbqlI0Q3sbUd4aFYnGjEBFRkc1gOO3Wr2s3L/VbB1iiqTRwsOjMD8rlge
2KeQB4TZQFgC7MIrlx2radIh5ffCa8Q3Cx0f9U8mA5e63WYnk15BkVdnROzK05yWUbWCoi0b1uVW
O13ReBB9qkWkDXl+Mv5K4uqPx+zt5OYdaCRfRcOlqXrZihI2FlJjWtZo3TEHM1Gzpp/gx3mC17eb
pzEL9DfTts3c11AXztRVsHmfkYjVYGCeIUbKs4DD8rTQa/KrPw/noR1iIbA1NpAWYICP63K4Sgk1
Z8X5biDe2R/V+XGCFHnFfG3+pzC0mCo8haZPfIxS4bmsBxDQAnYcpJuxjxTJUAgCj8O8yxU/Xfnd
/7BCyZhAGM6R9mqrpBl2RVgHhfSVVgCI4Tq3MZj/vG2aryFZna3ZLkOKwEoFmjWAp6zgAtwUjf49
zvMofrNbU+P1HA6h1/JYlg1w1zIUUOsr0Kdip5REvaTWFQ9xPUazjNIrb032hxfDJAQUNhApdKtu
xiFsceuMjAj6tXQUY8q4+Fe3ucf1gdwZpyJ3ImjXiVPmJ2Z0ozKKCzlEzSWLePVcSduDNZkEC186
g55OTElP8r4CIefwbdYsfElnpdAokWQPaD9nnyGprVziSQCAJ45WeBAnub0vGkPesNkriLLPgu3b
MYkVnzW/nuVsQk7r+HtclD8lPneoNFkiccw15hHCWDvrdmYF+qP0injsUzW5Ife70T5LxkzSrYXf
mT7MEzpGWUVJVxO6SGblp3Ftm8wD3cOp5mf91H1jRir6LAqyQSLNNRovqoTAvPSfF3JfX6llP95o
dHk4r7B7zEoC8GcMhVuUhqfaT5i+2/HeBRaxo1Ej7t5PfJUhX9sGtv5csjsAQxdUgYT8rKI6FQ/Q
RkXxCvlOoOQbkRxaYN6wmQtivgh5y9iwRpTJjQB+rJPKPmvuppbEMOFVI4P+SxyduV7IngQTiQFg
8kSg/J9TibQhmu3IhIp7AywnGcwt3QvNp03l74cF4t9nh5jpsH3dbxvDjlVqiDwfMsChUPLfAcES
FJN6APJPJlETwhz7nUodqwJk2xiTTKuGYZii2i0jEC/slJt5WS7idw3JAAHO+Hqf912mt9Ye/dWz
xCPsg2agGG03AEjP9p3d5/reZH2zmWIfyndKbYaqRVA5Mo8MBKFiAesLsSAAqm8Fq8Uvpxil8ZgB
6kLE0dQeepmJMRMlOciTcxWYKjxcuxNNwtCODDCBne7G28tRhYDq+6OFQMN24xHLKNDzgC7C986K
nTNnIXytvSyTNjSZden8b3PFcDxTUpQYy6Vd6VECr+4uQYWJL/N++dGHzcoi5q40uNXyKDOnsGpJ
UklfxeeL5uxr8A/1Q0N4I3BKsCb6mJFMjNksSTqTJy8QPNP0XJs0xZCIn2cUYSenHNRKYCltQPMR
XIjeykEg+tER8xq3iTrMHAOMv3lseDq+Pb9YOoY+1S3ASE65vqu96RTU3kD2y0u0W37HfT/+KaFk
sn9bo9wiEMQClrsy/z7B1nVr3udnr0xk9NKurNBy11Texk+1zwcO3sIgsgQ/gyt8g3LsVKyg9ZDq
T7KV8bGnjFAaoeBfmkzWRc7ZpJMLOk4ymdeRFvxfGmImgQJ4emcJ/hPlM5MVFJTX0PZ1Rrqf1OYV
fOavENaI6zK75jpWPApwWjX11hvyy8N9w6f3Yc0Mzm3ZvpR+CV3Mu6kk0nGFiUVntWXNhDbqqOSE
OCA6cjr8PaS8hx03XnQx3VFsFkJPv/E1d5QLUG/X41bCxYJ56VeilFmawxVq23UyGSfUZULNrEwQ
9enmtD3VWPRqXgIUGe5rTAMLQGcrkkIHFORefbE9WQvFYEJiauXi8kreU1/5lM2N5hZR51bT0DgK
sIqWNrWMFrM7sbJK64LQf+4BRlCvhREI4z1mSyMo5b32XZKaWKdlBHLv6TdlqRu/E2UrkKN6H/H5
Kwm014LQXCzyiP7/aGVpt6mX4ZfXgMsGaDltxOtfy4ayuAeIrWnVHQWBD6YdJsufpmxw59BxcwCq
0gPcck9dGxkfEp1by9LTp7vN7llqaz/Ykw/Rnp+OzDjaXjr33nMPWCwxIq7eiOVQ1gB0RgAJs7Ts
j5rGEzwjIwC3y134ykchGB3v/eGhKVkVC+b9dqQYoUpwx4UWy16ObWR+f7TBjF1iM1mgxCqGD6DV
Ab3g3zNbYzYGOT1ipUXkKfWCu1Pi01HW/kOSK7H7AeEN6KuJz3zEiYlsCUg09F/Ptbq/lX1rOY7H
70vtDcx+q71QAOZlC2/4+u73hT9BabmMn658/KF32++KwQ+iunJPXZNVr2t2DkP2Tmp9HxyrJXoL
++VkGLSyxoRz2UyyRq0eeViqYoU+DNaCL2Ur//Y9g+JAj3eHkIRLmQ2q4H/g2d4PyT0KCJLmm3dj
PxDb+Dt0luX0j7FBnYjY7XrjqPLXyG+7+3uanxrccVjXUEXRVqSz2xnu93hUyGjhjr8zQ/+E9uAz
daqFssz3Yx5q06D9E0v2fuyYWQM6HxvSwPcriOi6dptj4+x1QVVKT31iM8aiCBm16oCHfynZIvbL
7SWV96mQrzFNwG4tffjFXtEEVswPE4JALWY96HVV5rtm3nSY5d6jgiU6AKyQaTj7i637WiR6B72g
d/NVBu/s6Ha7j+q5CWpnEEG4wccVddwPr/Wzzhf4X4hOeUhzbZCvfvz1J7sO3lbjyWMZl6cXxUex
RzcCP22VDWZTgrqOGzt/w/OcpYflfHRC4uqLuHkbZtj1x+89bBFNUJiQzmZ1G5ZxX55myUdsn52m
zydPOZrLrS0XJDmiUEAS4Onox6N4jlPMkBeGY6swZZJx+EZP4EW4F7YO1Zn/IxGG9BQBIDYbTDbe
mOGvcsz0l7JQzwiD9crmAqDQtcELw8L4DsoV0uD7K+PYstJ9bQpnuU2QWmHSgE/6+b4ts7/uqwRN
qvtQfo/zRLQ8eQJHuCcX80EaPxYjAtMXgX8A3c2t9FDch+/acywnBqAYhUmLxzedyVpQ8KlRykeI
7XWq3ZoiESdhEePnWgQtdPQHs6EiVDIVVuL7/u26/FhHoEVqTXMOmWwMEX45uxZTzLgfMajK1Kjz
YgjnbJPTZi2IJwABzWWhHSnj3X5GZn1hF22Pzz5TnBGLT/f2sbMVBVB/MFYVmR9XpLCGMqdEtEx+
OW5IsyqBFKEyalKWx7eRCT/wF/uTCK6Io5jI9vunIrvLBaMAXltTajMwZfN/R/Kvfjj970FfjYlH
0Dp4QaD6YWgbMEzxQLvRCtweu7wBU0XrDES0OlOxmL5MH1rtqKEtUfM8djYMVWH+f4yXe+vlTPA3
JAAMzG4E4gARlQM1Ds2YvaZmxsfeDeZfpX00F70cMvdC5rjeFfzYOlsOqO4XT6idUPmmumebQ9Sl
DMi98EU51M1H5Gs6ABsJu8K9HBWyx5sfvhZ+/3sBe3wo4MQG8MVF6YafMTSwJphyUjKIYAsRG66v
KhsAC5B3RrHWJHcuNUk0AvPlbCUeiTJ8k56NfC+dVZIGCo18578+Cv2n6hFn/EfvBQardp8Q1d3K
eBogFJLk+NdE7+KrAuqhxLcrrXfyUXwbaXKzJM2IKOg1pvj6poRZacbVfoT1Wk7GS8izVfqYSAZL
M09WDSXP0om/nW/yodcriDHHgl3HwCc8JxD94NMREJf9Mi6NnLfK229S2egX04r0xxPTcfu5GEuj
hfWH5ahflZMfAhB9xaa3UziyEHUVeAtycAEZtcZqqAjetvvH9L59jiDRuVMu1wU9ngrxq/BrnMAI
1ZgVP6n3Pm6noltGzDvoVWFRFfaqF7vmT0Wru1sFQb80wKsWM5UfnV7Jb+UwRNe3F266aVbesZZh
hBwkvi5n/7dJNIp2MI/UGTo6mVORewl68WCbtXypRGRI4b7CWDeBrc7FEA4ik6QgaCtKbEHivHkP
SjvqwBuuWpTB9+kLeqjjuRy6nYrMjJbFIbBcKFkrsAO4e/diow5IoLeyqsrM8y154560MKfr/tCU
mHYh44dYZtVxsfTkU24D5m5L/Ao9ZBuS0wgcXibQMk/JHkIF0KgnASbQ2e6yJDuJr0LKc1L3F1Ji
FJzurlUkLMlccFX3qLmI3RinwjdBPyeFaOIiiv88FKseL1tsumEX2VFNCHVHlQLU+8ZkExO27k3U
Xj3RLcRdItN65kEe5mdF1hpaCwWi6OpkA4Obt2q90KA2gERxKgWJ2v+i1jz+10DI5fvBtMUAeQWj
JBBtbtExG3FCNLPjahwk7JbavYLcIh0GinGoM3oJFgMQUQTGfyanSSSj5u4H5/pa84AI+2517KMr
PSKdwoSXW0WnETlDroEGb7SlIYLP5IB8VhagGmWRYSU/6HQvwt7Y5z0+Wz4v2C9ZrJkdNsrOckPN
5IrVCQExfFXZpYAS/qYT4yaknuLtBxVqrdLzVLLMFF2ijUOEcXrsMDv1B2G0iptCmlNewTmSGme6
ZmBV1Ymn0QS3nDBbyy6uBs2JhT2jMkmYo0Nl4REYhn4gv5itTablwaEJUuKEIM3am5PosGRUfU0x
X3eswqJ3VVXjarN6a2F8+42ICDqneey0LzvSzJyRoBWsVssrOBX5KKkR9BL3KEme2ZolQdu2NwfN
Gp8OokvVg2clrdUTaIDa0qEJe7QoLuWZmOwGCe2YgUttw/QpS3aLaju72P3z9iGjfDOsbxgpnhqQ
MIB2Mmy7iEzYA+BMPwaXXtSN5BU5YWbOjjFCIAlOKCQKWuDEKzIYZww4R71c609/l/6+Jo4dEBDg
u3Id5Bvu03CkYWMw5JMn6x1MS1Rqdvw4+ObSFVSN/flcrRXXX7B+eguTPelipNZKD2MzILnAV2aW
GejRGGD0E328YfBthjq0IdSyTi9O+N1E6pJkTZoAm8QJM7hi6Af+iwavCP9P2UfukcJy9a+Lw19c
0ctpL3ls3iRdYWoMKGuVcaKjwIBEpcCI5OQDx1VMFTmry00OPueif9SDNNJAdk7r0PDSyaWPat0C
azjsmJUAhhmxdz/9Q3wTTuiF8LbvTptyn+doGhjiniZMJyrvAsEvkFL4DEZi4YhqjirnKHsteQij
cXedKhGPvAe7HcfFxc5CWFbX0T2aYodfaLgzviw+tmPNVJzyPLuMPac9wGqGK8UwiWUfCYpQW3Q9
8KrDJn/YZqZeKH2qJrDhyrmYQz8beeoNGgKBPPhJnHSiDuXPLQ+KOmbP0fG1hpkhwxJTCf3CbjYJ
nJFbP8jl2KjLjg8i/ZORwTYEseuF2Qxy4W3to8vnASEiV0H2PDGoM3gUJ9qvjkpYD+waMFQ1UUEz
vGrf78f5aldinlvH+shqa6IeWPu/w59kZeq+qy9ipd9tNC4hf21Rqrn6BwNiH3k9jGBgsXVxH5XW
IegO15M3gr0np0Xqrtlwngq5vhtk5nycmtTqQWGII3l4xs+/a/I/X3Phy9k9UglIinLeYCp9CL8Z
2QS9ugyXLwaOqwJWk1FpUDPQ0h/oWzJ2QWDMK/JSvF1l1gagFykshh/pPTc6Ccg7SdbjxQTBx6Zi
jWBG4qGB63zO15wb5R2Y8ldsPTs7lLbrjQW5i8+4SaJRvAPGuGXV+SfhsLcSgLW7E5Kpqkud+wsf
YSW/EU4CHBmHf0f5z6uvZM5Q9GC0DMfzQYQN+ADDVs8OV7/3GI3/AAaBgXtumktuNdmBR/GVXEGq
MlyjVHvfMdDOqSu0WO5Z5QD6mlEnkwLBn4EuIJzVt1ladg2RgOwbkojUiiYQ3ONOau8i01t11m3H
oITKdSfA+X4UUZ/8Mw0ZU6HZPlmBTdr2nk+lrWFjetVUFYJhZ5n5xNf/KqV5es1jO8Hy6UGrNDhH
lvaEF9wdrhtKzP/cv1uw5vU2/COcEwfTjK1nLA3fLd4zxyMWbVD/F4ycGns8eFcChiqdH36nQRuO
Y/cXdUVhQi88HnZjdfjrTzVxaV80SLmGYw7G+SED1ZFlLaYQAT52DOcCl2eex9NHRpK4Ck1KNJNS
BTfkjPtt0IIBVjoj6l4/TwZuxf/NoIM1lLUc1vhMXOpWKsX6jrXYa5cmx8Oki6xkQ1EhUBD7nMd7
zNGixLP5FWM0Mk84mH1NdLhK76EvUpp3niGc/z2y7VLhRjwZp/CYH38rMdyKsYZiQ+b7/ajEAcyt
gRUIGMPyz770Eplea6pQ72ZnCsb7JPwG+LQgMOsNogceTTw5zKxsixN/vq8gyqsvvkHS2IVRZouu
naxO9+heRvpmfCbJkw/f1HEHs3KZ2nXVv67dRnCaUEEwKBsXZcJ8C/E7DzMxJdL8X0ZOs3iBJSuR
lc6ugALncUr0foi26Ax2GILD82bnVoaNcG/Z0LtcbMAbGC19r0rqvoXS+eVE6shAcWvHZBPLJStA
hY8HpGA03bu/lGpfmKjiiTHXKTEbCSu4VNYVS7dFNPnTie3eI9JpKHxPwGOJxDy2EAH1yrDa3/cp
H+0E/PwsGtLP4izpDALYtuGC7N2+mu22VrnDd7kN7UzTwRLZvKoas9iKXINdPAkOKvGwqZ7Fk0vO
/hYRrqIKX5Keylv0D9zh81qbGkVYvCOkfPtcpE4BRQGuHOFWbgB+r2JaERpdYv4Qb67uGLGxk8MY
ouv2nW9/Bbs2dhuV2hOtf9UzEdbrBCN++LBtuB0VEIGsME5i49t/rZaw2tqQfSO0pw7x1bGbv52g
sss8Rue/Qr303uQkbapi0W0ycxzkrUQ8Uk3qMCO5FYjxjGvdJao4bPN6+qgSHPF5/j09jae4g9tj
DUivxkNnHo4pOhkGecJM/WRBk4Bo0Q+VtRRjblCLzl+0/UdYQrnz48rp9xaILDuBjlY4gWduFhaw
WwVHHQi2u4fSarn3U3ccBI8rpp/6tzvCRMco014eolyHBZPv2RrcpZbT18jEb3YaBTBQRKBfs5KQ
YQSB0JqMVk2WeOf4Fi4fEPhEV7X116Hzg+EIHqxH3nWdFdF5nCsVgKjzjsVW50bfoDsrcx/EWxm4
C8vDNXLl/QQpEkZogdvXevuKD8lMkhj6vkNMLeOuHXtVonKLOlZ+4fi3zo0ehjRXduIF42G5Z9Tt
WRjn0JoOh3+oXqpGNeYUK6mfzdCV0HqudMMJ4tjYJQg419jL5ZWt0NVUFyrXTviFrmglgDy4Rf86
5MJglOrGh9sBbB2ZWo3GM8v5WKiArqVpxBlCZshlebDRTHKSWJRLPIxliILcyjVzdsMrQmyaJXqI
k6d9IgXGlp4sxCVQBLUQpw35qE/txiwv+D+70/l7k4ACQyK2eI2KSsRgXePMx8yzaAiZKh1gAzgE
4gcsT3aLn4iy/qMyD1z4sw2flp/ATUkYrymiTex9b9sKG54pDP4+CtLxplJ+4aAlQP5CYnncGYrh
BUqHd//oexT+GXE7+2FPalkN6XnPEPF9PKY8LMZoiCpEnWtJBBouGBYMbUp2eV5Tm3EaAHh6gSrI
mBBFBUI41az2lto5BTWbj0vmbbuoPn8WEXTVwhezpf/eFHScBfAKtEeGs3aggrBSbnkwyKPW1f+b
A+fjZEkS9Zz3oIVhWrx8Kd2mdqNbQP7TThGA7gaLTtFbeSzm9p8zWzAE2hR8A2qGhwIInuMqL3Bw
Vefn6Cj9eWNwkHVHI+BIr3XNfdn6pdj8tHNE20z6wwdDiRzj86ch9qTc+CkSlZyQGOFQDJYkCwDa
ni+CQbMazwUtupqL9xehd3QoPUdyVOw6lEXAIrMJNk1/D1q7qY0Rfh7XzMPKlnNZJd5nexusqliw
kErRjVozBr7Iu7126NkMuyNLXw78MpyMAm/ckyc+Xf/ifHLXQP2dmour8Ou+ed+BsSxO1JNOtAl3
zsMOAA4d3UhojN3ZfW2weisQWt4xU3vxIkbmE/nAcjRPsQMMWPzkbnH22i+srjnEdko0wqtlV4rn
cq8WyUwNNzh5YTo0EutbAeFc4kuyA0pV8EtllPaOI+N88Pf3zR7IGpfK0rVliNbUQIm6HJYbYubH
hkuKaIo4QeJs7IAAEUQ7xFCcecG99X3ctRq35g/sKMy99KItdkcMFK8zgF18SQ8v4ktDM+Qmv6gp
oPsVcGvwqQJzuU5EWRKyaohvfOhy32aH/4xMnEoLdfSFmlUFset5ea/MCCSpVejZgzNpAxDTolUZ
uDA0Ixr5tPeX967QkDvR3bJZ8hnes0FvWGkl8xBQnFtNzj132KmfSY5TgbVyBtgSZKonwdwk2OnX
7Ew8YZbhHu/RIOHrHMixL8nL0eooTruVCqUcGKza6MVyQutBm/FS0DMjvEGS8IrZRkn5528vunpQ
3PbRprD5WK12nx4I7N/PX+1ZFONBiS0fhHX4rIA25Y3mItovpmy3ZCZB4nP9cLCUjWDY2n+hz0AT
gA5r5Sze/aOnmk82S848CYEN8Jh1+JL/Prm+n9C4qZKkTYSkXiuZj/oPKxH+Q/EgrA/FFkQzq6e7
T4/T32oB8IdZ9A8+3EDYqeEtnHA1KybgM4usMav4QqAPUhLJV4x6OqpJfdHIpKRmMuq+PKptj8O9
JHE6RKYwdc9DRnZd17FSouWBPY5GoCbTOozxPNYZqaurRtO35skiVrUsrti9/RW6VQIwmh93YfVV
CPbiLzCfJhyXPLO5i/sQ7tYKyIJVyDD4og59aCSbFuGD60vVUDwpFk6mfkJtmsDX420qIVOxyfwU
qFitIaeWy/GQMq/HgGI4HQjIfc7XucrDTobDt9qqBMRcfGpksTr1eha177gl8s+bJCTZa0FfE+3k
UzYIw6TxqjYzWDf8ixTlC//+xf9yolp3i9FrNcmHBDA3k9La3YsTHkme0XP6xenPXqkF6avd7AiU
jQ31H/OKaEPI3IOAYuVJyC6TFPYQ4chqZAR5TJdtiSPZsPK1YjY/JUOPN17Af3/l1hshdpvFLdo8
a6+9tHVzxOPBMwNMED37RhWvSX6V9y6eh81G4mWaH224OwDoA4RrLYGgR5XZhcb5UP+tfukzwPou
PpKKYXJ5AqqnNs/Q8lwyWnUIkO6e2VLMvUUSbAB6obyHPr1sDokC7MqxHNBP7OXRapK6RfujGX3+
hrp5LHU8s6wpvL0KiGIGPMaIu9qG59MuhDxcbsPaQXXTjoJWl6jKSdLO8aJ4EpjuSIXvb136LBrb
uECNRFJTncyHs3DLbq3qBKAI3UXuc3klWUQUrprJjbOrMDUb7luiQ2jrWricwgMms4VeNeTZKYS1
kwPSaH7m6D8/ref0/5dqu0+/4m7PANfBtGC4NVmQPFk6q+Mhj2fkCjRApc/F+4Qm4M7GeUlJHSno
y96aUwLj5ne24x9ZodUXo9HpTKrCsoW0hbVhl8ZrBE45Dx30sxrbI9xZoCe9Xdy52o2DY4NJJpKH
ofseBIDKmiDamvyZjWcYk/n2gpEjpLS4xTWPgt17TD+oqsrlbKFt57i+amCoTcwXYLgJwMcWwrmY
efugmtWAHx6SpLYl/d+0y27xnuhMt8OCcLxubW6qFzmEtvZIPuIKJMuJXX1HYVYGGKloIRRwWGUn
jtQFQaPaCnDGa1MqhASiAL+p76PGGSfALqPyYWJkrr+SF6S12oIdGnZV0N1t9iHlWKNXXj9NPlt5
RghnwZ+XF86fnLi1Xsi9j8aTYynJr/GJssTPNJQwZxpmh52fAFOjraV83mVhm/5pufB/R5oNCLqB
bUFZE6n31CtCzRp/n4J2pHAj7R/hj70wviLLENdISeeQxX6ebE0Vs7JBCAktJ/K/pWMf9Vl6WgYV
8xSzjaD6lBNeiupz/oDHYC4XwSr0NAbibm3p1OwRAnEzKZvtqDFgPrd81z4ESS/V1QAqnFOdY6bo
GGqmVA2JTMuQj2j0vCxjrbGh7yFwnYblXUMa9+c00iY5zrkzXb8Gf8kim5BbaLU6SZNjJLPM6++p
zlaNUiHs2z+xcn6Fui0KMunIVnYHsvpo1L0lP2vpJ2+KpbWchrZJ00R5SVlchaX9TGv1C+UaVAea
K3iL2gtKjuZe9oBlA7r9pwEllgyxz9MBiI51dXHBNoOPyzNtAE3MN4zmxmhESo4PkP2rRj3tHVUG
Jk0aEGad3R5iFymTTID3lCDTXV1WVMBGoodQNKBzALozaN+qMn3kB3hAggryJr26GK2RYYLbl+Ba
QNP8DsURw0Z87gpkAU6BDsOfvRr1vEfjYtHB8a86uZa2S3hV7h5UlsU/p1LfK+/F1Dlxi9TdtBew
pKLAgjIu+fSl1aePpHQVd34N8CNfZBxx8Kuej4sZLB0ra+gCdXoeg0lrbl2vv5Y4pJOZeC2ECF7C
t8tDHE2F6qBLwfU+BQvhYzLBa6fszW8YwfSd6R2p7W/bgr6Is8aKMOG12JKa9O8WnDvehlGueA9P
55FaUBf4nw4ciGEWuuTwcqiTAGIA2lM5lgiyq3fopsDtStBySMhW355DFlIalcm5MzDoVPHdkhQD
KJayyywn6fkh096dmkQw0HQpUoQVXNsziHAZg0lg0jdahIDPeuDlf0+KFSVxfLbco9Uksnjo/uq7
CzGD6pcyzpTb9wzB6wiO6MhvnmgIRqKao/OVuwlLHrppEx5UyBn4b1tvIgY1LDUoxhjGIlKaJBGK
dOt4d3giZ1p1BLEEgQ4E4O+7VVlTCY4coOton4i0CrwdSYE1ablgVA9LwY/ItbB/gfM/w6sP8Eu4
0lM65lvs9RvRKyeOFMWRu0OHvBb3c0mTDuUMsHd7wgvkNGF2B3UTyi7q+/kXbRdODAfCXMU7A/El
t1vYCfn5dsAL8+nSp3Oy9WRX0Ck8nGm04yf3D9O49uC2Q7ruFzoc2NaKfiqZOE3ErjvWwHDm2t2S
fLCN0jypIYViFf0DIOsN0P4+TKFJ+fQmRNoJaGgvx1te0q9nySt6/QZIMlPmvP4DfWOFradks04Z
b/DRBrVkRD36yBE6RdFVvIG7NcpCg38wwrX7KyAaI6DczbFJbpe795EjGtbnwEmlOwHvrzSiRK2L
5U0fMHf63W8cTPpNOJbCG3w5tWI/nLSK8i38mM45zxCAOP+AeqWQxSxv4XWiX5ai7IMZfZG3Ef5c
WFnTZYTIvjpyJKt1PQYLfJRtZikHMQYSNd0tb4W8P+oYx/C5vtZucYou/eW67aMiouOuxCbqg5hP
4syDDZmkDqUhFAQbo5V8yZRtmP7ftljnbDyZmnZTcyfyVbfyG95YRGn4ekWiixviIuUcth2AkNGA
uQjOvvFoseYNeJuJ6HiZ3oj4F4TF/z/GUmv7WnfuhzzdERf28kgx3mDDinyGOLIGSNR/jHBZROlu
DgVwGp1HX5NNCrqCD4CZa06yKe0JZB4XAPfGebp02JdJTXP08x2NYKMxqVb3ZQQMe81YF+0Ajh96
CQweGRfsSZlIkYIYV5GtqchDF4zq+RiqjqGxGEWlJk3/ve5ffQFePNNLjpfDA3cd7Iizrg+XhRLz
9d50ymwgFfujUm8pFqRES3aEcwDgTpZaYYRFlplKo1elafdrrGjtVj+aymilI9u9i7oB10TFIxy6
/nH3br1IWyZsPRSgrX9nVWkuLkS/EiqixOFZHtIP9B55F8+0QKmNV7uzhSgEFsFGaGJI92nSyKOC
Fb0sm6Kcq8ZFQNr9Kou1LD1WhZMP1OKaD13u5YRWLJf/l6DMvfReDT0yyMmmIC2/7fL8ezcYP3Xh
QdL1toMw3GW7XLD5v8KLAJaOnD7Asgmt3nSoej8p6EAqRwwP8BB5Icna8jpT/zxhvueyVdpDObQD
mRRGgE9ERQm4SuvuvpNxc+t+tnAWY8KjyfYRwhiir/u0obRMWTFfYZArBMsQesIdH0FKTcfeKj4B
Mx5yCq1eLNXN/y+SuCWbaBRWM6soqX81KKBlg+oxfA+3Lfe8VqQlP7+PSztUaQ1o5oK+USrY2kGp
qYdgt8SP5swkKP/V94Ph3yfFvrJKcxUNL0SYqkRuNquojBho77DvWGws/jZrby9Rtn5Kjq1WsJoU
bs24G17Yuruiwc/o0lxwI6O3FYo7S7CZ3Le+kRSOe+prgVk+m2TH83n7o7J7gzCBOXnqW9ZFbjwG
YR05NLwVMSBY0EBPBmqSu61ddwCe+mYAXbGl89d7iSZPh4qHZuSxTxGUjJwk9GlcE6OzuuWrjEub
8GEjsGbMNrqVipZ4jj+QBgojhSLsIc/4c2y0k7CYxqyGBwXCvAFyLZfU9v4lOoUYho0qiotp9wP6
+Qpl/mI3i+s7XmrHt3GCo+q6v4tywMY+q4KL569+nX1zkzdR/4qOjapKtlc5JaV4snLuL2VrPqfP
m2Ck5kbucPIHymFxVeUJggTS33xrUrssyVjxvZiuUklxu+psyxIt1StVPvpzCHwXUQiaktkM7Qc+
8knSIjVjgbC8kOuYNH72wTmYGrKg0NQxRhFTFL0kwe3tWpeB03Neu8eNxiaKOmLBvAdc0dDjJX87
zFJxVRvdCuOT7fzokiNRU7ArTTLuuNXqO9dhNR8rnvyzU4P/P3CaNUofJjWJ/0CUsIvOrlCaEwfz
L9OWpGgF7NfMJ71HpXxFHb0gyZYKXBLdJhRsADHIDR4CuS39LuVaBjOtFbPLpM+mctEoIVYBMyPo
byzcF+k+qYxgv8OwP6dFrQfQyR+mBwxjfDHSTqliuKJYZxo/x9HLqtXhR8w+pzfnUwPG2RjJL4R1
FCILkOVOPYlb1FOaPiLzKBDi0mng8ao52sDE6aud1Reg/OPxmJXZBPsCFD0DYFtSC1rO+hbeFEUe
ZIjQ5w6wwLQC1E/SCsHh6GggjYYc9x9wmA8uhk1MymJszL3xSi918+DbpbU8p0qBnWHBeVSOGs8l
HzHB6cbUzDwy/57K1e41XDyyZJJ3qQR5NqLOh3R1R9XYX4/87CfA/98ZdeQB2YP2EtskySb6NsUh
DXqVTHGP6J7aytoyDnQNQeo7bcdXekfrpbl/CmeBIGZotYizkdcPpYdj5RwNyJtDWaigzKHyla6E
JpvNqzei55mPBj+JA/Fsf4yA13VAfg/o336GR2gjvkgDARlE4HzBxYJxuiN+7vpiGd0nYf2rR3V4
PX8u9snVp28Jebl/c26FvG4D9ASnD2oCptip0542dAX/ronlRLY+3nfqXRVwffUpiwzptkUmqegs
XqxCMI07EJI/XGu0wu0FOaOR3xxqe+m7wPBwLWthDgOdUloVbvwvyZrEITzNBy2UKpM/OvTmPJCs
ernWvRuvspDiHlfy3toL/vgMTGKEcZ9lI4Gp6Z7A1rz+7r5Z6E0Qc0Raxq1GmEsbn5MuiwZQx890
eT1lgAgFDzhA0W8FUey9rIxaPCps4TcfApSzQP6zGFeeQW3WMo3+ssHlrWbCoZIKwQW48KGRhdlF
Bo/NTBlZS9CzycgKzybMvCgqz0647oEJrcIsHUGj/qp4kCU/+qj9/VYQZ2YoWZnOx1h/xE+cWm1W
ELXbT/6SgUZVB1b4Yymg2p1HkDJwBVw/QHOF+jlpCZ1baiq+gL7J9Osj4sxiljHu4zuPHvbQdeb8
e0zJIis/emGRVkl7KWnpFDgjRblK+sgyOl/YhI6wBh7BkSjae2hCCllf9HSJkbsN/N8ozUD3RkEr
Xwp56YJww49hmSo7kWNPfZQOKEj6yu3IYqkAGbI4aFnAyxLgq+3sZsxcK5aOmkXZzHBG742zBuCm
BoponY1FnnOedk8906Yh2AipzEQ1UpgitLPZeaFd2R+IG8uaEf/wWdzdTBu5iZXTY0hCnpQPRcaZ
lXK4gv/hjWJxQIs88hhq6fnAXV7eX91lr/X6fivfYbXN+Pe/Rxp44w2OCoN6QLxxM0VOuSqAuwds
vfWKozx6M/6rFEbzlxt2D8T23BS4TpWUcdAlEGcepb6sBf2/5fwGr0cSckhnAhTdgg1x36XVYnnJ
vFsFSvx95jBCOdZDhDj+mz61R75wxw9i7ODo+iAM5U2O+OyHOP9lYyqmOCkkHpT+UOGtRf/lebfd
G+W8C44WNCJyFKpVSQKs1bFho21kVTYqtfXTDZLHtLBo47aMra6zqmjzKyquQ7A3EXxlO40LZDwX
3CF/UCq63oAwvMGf3ehHt9DIawi0WcX04HpZmQxU3QxJpC7UPjU/8SRoXUC0/d1994dc6pqt4n1P
lpieclDI1WyMdH9jYoi+Nq/jXiypJJm9ABmJqdOXeUPixoVRGZVlPnGjykKMjnI/sUuWNQrvoWlV
n5YRaMApn0WhxTI/dVOh9cY5c02ECO+oR+8IwxpXWF2cnN8v8FGEFvRuQF8DnS021zYzf6UBX3iV
+y8sEA9E4n9YcPN9EDoGBDCHOwWj0H7dSoG21A5PD7Mz66OycS6c95fYRQtEzwkc17uP2W/BJqP6
aS7vilt3PCh140m3zjYnjXmt21ruwr1CibF6FnMHZ4mYJt3pVeBnePZOlwcPo50CMmulYZ7a0wRh
iO3e9eX4eJilHTqOZ+20xo8gvXO+dit3YTHizgEyA14ZSmreyRI9cw2yRrCfNgkcp/U4fNCPCvx/
/9v/0Usy7MzI6WFkb/t52mnHtLqqOQZ2AGJmrETcRLkKaA2F/Guo4xsNsRNOipwxrztcsbXybavu
TB1cL0XOdkJJvR9z3k78+H/YmytzeRnkd3inCydW5jJIwzvAUDWc8etLkGDSBQUpzYN15IVgOFw0
Bc6YBk0GHV4L9f8bKWTUKgQdRG2jT21Akun9cI9z8gGn9gGAbmnQjfvF5It0zMkqfqck6l2NOqyU
MWz0hY7qt3aQED6l+/tHdhi5GDWfarN1gamRepzeaWZCrLGxKSJNJK25PMIrKxoGYN+Yb/3JA4YY
e9yC5/mUVgfEWxjs3bdMdR7D6COCHoFh+WuHHPjpTQYMd4cMMJ9e0+OnBynEK8QCl/hJusbllv4k
CDdrGPhsZAuQPJ8DWnPFZVabIDVERMeyCoDIB3hpFYV49WC4DdElHFRzQnWCQCFBWLhIwXS9Ow3o
l/LuQbu8q1xvHSWQ6T68ClhSiFeRsd4ZDXR2X1qcbgoyYe4ab20p7ICjjwZFd6YhEsdtEINe/AV2
kAucoJxKDcuQJPihZeFlABE6/9Cke7tJ/DQYt03WtzY/2ambxVAjwm/n2WbWLBTaazKeNvz1njUM
2ViYcFRnEu17VcIdTkqC7kRRxOtqOybYCZ+cxiyzEChzlTkbJkp3atCb9ujjjGSuy71PJtUv8AVR
5J5BdVRAhHOWjnzOIeRyhQhGPP6iMPB0VwfSalyn8EN8qEzEMQvAcH/liWkLQUrwEeV+RSf+ORz9
giarNVWxLr0liO7gAVqmo04KC87kAyzz4xOFzNfyBnWErXrDT/1IIzolBbdkT6LRakaPYl4UP83t
eNk4BsBYa5Kja3dQ/6HDjjV/meQyjZkLQnXj/cqd7Mh6Ul0MntWsxd301Oh1FrcHOlhAS7Pz5+Lu
4k2X3SteP+GGUU/2pby8mZROd+D0v37Ulimp2Be6nxVprZeKqoXguc3YD+aGlCWwgLlvNtoEyXWT
pnYs3MjBnhFL7yUp3/eVzzaIm8khGM8t8TTmlc+Jqk61QumPOjqreoyYXeMNzBXEdwhxT3D+aobF
doMVd2qxvtu4n/tApE5uRKdF75eBKknb91CLjdwJVEhsA0cx63bmiteq1nZ3uik1nWf76uZBpw3C
yz89jEaPqu+TXVyfbYJS9byDTOiXqxUGs5y8HvZNhL5N0+qd17uBervIO+ENRqIOkLXKgQcHRhRV
EsSGfYUPHoq0KKJQbtBKqv6YtYkUyrkajkzESJwF//K/Lsrm+1OkgVS1db8+3Ex50GhU6hGu8kEZ
dozoT2IVjqRHf0GkTqPcqJiUFVof45dk5n+VPyY12LJGZItJW7oEndDdIYkwj+Pk4vnGUGmAkiCB
c7vtQE0fA7EeILvm/NakjCifY9UCPKcNDOie4RZ3tDSe+kj3AbiqbHI+p4RDVyGjjhy8zZp45knE
LznmobeMtY0OSCqquu+pjNKEqcC60B3h2/FwmyuqgbUzPjaomDUYooKiTZBquZGABe1nNm5CI4HO
ODDW4QAb+GznuBDeZekZ/mo2Pyw0vZXHLIurtEO3jWCNLdHk5tuUrTF20eS1QExfJj2dq5pLt4MN
YA1IDSOEKfYSqSdQxvCGO2GvZ+l8txzoTnuurXeaDEv5KAf+9UPJlBZxfrJ0+y9depfvHhkSuH3g
Y7PtSqDcTr1SumgO1wJHaqVKeR32mPTwRpWgmbn+Gfv6F9fILSGjs8RVdSA7JjyfJcRYhTuCWVO0
GhTgG8qoBcKHEfpxIVVoopprQUkS1YWAzwDJHC1N3Xm0TrljlsxVHpedbuqjREpHlsx+gf5xSv38
dNAN4BJK2UURJCEL6pSK9q74DeDQJuv1cOhNRNTeW4yjRYSesNELuX3wnW+q523gokv1NExi56Xl
/OguLQI7Ih+dH+AFMI4jquZkdz5EJRN/xcWBmfs8aa6JiPUrvSjDCPXp4GZuEEN25pyj9FI0OCa8
hRLQGfczil5h6ZG3BjnHH7nev+xfcir8tyM2HQDohPGZJN7jTjtnRzpZO5hZfN+sEoF4c7F4p7PS
Z5E7sUKDQLwsdmmx789OMATNNxoXjbksYS1rfoa32Y61o/o6pUs3W2mMKCUbAE6kFMn7k+orcatH
AxbzLxlQTDCoq+5ulghn4ybbwakfIeD1ozRg3hCfMX7dQ6SiJpM3EQcfUGu4xV7GrDyK+hGX0NZC
KXeHn6uj2BQ9MPxHDHzEZGRx57mjr46h6Ur2xpguIYVGlcMT2804LNoMAiCg2/NN8WlJn5CmMNfw
vamA/CHGwu6WEtOXRjXWwlV8J3PeA5UzXz2XsjdcqWKy9/czjX1cD4adpoOsND4IfvG1XdHjN8Gi
ROsx+9RI9akaAK0cjaBvnxwx/tipXTaD6jYFzgt9VbH0NH90d//gBbBWxm3u/40Ey8SSR1P0HSc3
z2qkIHZ35yvzzDsdVW8t6MHgnIvia5chPOq1L2/5JO4yaR9AJlhjeJRjz4Ej/6/dvU6iaKdLcb4n
HB6e4J/uPAFFe2r5qcpBJoKhBgOK2pidY3puB/6IR75vkClHOozubgjMQKzcwu7HFhyAVdR4t3Rv
NvylikOmjCAuNWWLuxDBwQ1niMNiPP0XSrV0TWViLGxsJJ31F7bw//sZ6o0eM7vOXo2658OpHHyS
j0wGjOE2fNEGDXjdujZHhV4nwBgTrOIVh8xaLj1rlTvoTbPZTYwe/iU+JZt9oypM4PLabHUz5kdY
fZEQaOHPq/hb+nvzEVW2odddMSsLPfDqrPIMucIYuGjNSPDS13N0w44klQQh6qmHX5IXAf4gsjJ0
CfyEypgrK1KBrkCAsiVwhhYX8+axPU6x4rnc2/+guH6k6b2Mmp+pStLMc8opY69IkAdhmafzf7Gq
zLum14qrgvIf33vJN1GN9xCY3yMXCso4GGZJl6auNecUE/0ZXI0GfMNfrP5MkXEWCttHlHYjWxWZ
pnQvgFNwaxOU6iLJewooMpq6PCyQi65Uixe1Iy81kRrkQ9BXzYDnmQJSfIyWQxPePXLeLStKVNU+
zspd6UJsmUFMmUUqUzT+qhn+hZuUVtHAKwsOu/6AEx73AaMmbTQmtIHQ1fGel+TMkscAL1ceFIGb
heLeDkFCrvNraTatWzXbecO8xX67F0COGISL3hGXEDDLp6r1Ln4aU19cIfX0arfLF+HWtWiYGAT1
AZPpbUys3aG/NdWN8Nims7VbRi7R5Pm6+rudFI1T8iZWB7b5vd9g6FtbWl+prSPCZ7p+/jktYuca
qNHPu5D7aZ3PDqgSfNtO2L+wet5wJLE7fsuHhPaVHhgzcnitZxbu1Fl3IJ/FX9M3nmJ7fccp44iI
Q35lUSjaSvcN+CKwnzq0crbuB3MA/OFEPqzusw2yx50nqLFQwIl5zE02Ng8Fy8cdybpfixVexJnx
bzv8VlZMdQjZZAJEP8/JDscvn/VT8MOaE5C/Ivbpdsc/c7qth/2Qz584OF1aZQt17Btp1v2foVVL
xiGl6KDXQ36VdnxgwRAG40YcPAnJNoO3IPO6AFlAC9YqsgyOQsoQhRMKvCJ4iylU1NmMAx6WeFF4
BwB7cPZxWR2iyazukJXM2cKuEvwPbYLT0KKnc7hDPBRMeberKALigCk9wSK7Rd1JxZ+4UZEjLO0t
2LK+WeopZCPrD/JcSClnAEqkT3gQK0xRSueSsR1QDWQqaKPwihrRYSnoyIUZp3kYNZaHL9aZdcKV
ax4FUJHfKGBz2FhAGXbP2MUsxSItCDWVfOejtEvOByUHdMtEe2/d1m5RnIAfqQ/I1f42aqjj+9mD
+pYXQvH+zjjV1ZdeS9NKM1Wu1wF9MG/OCno18Q1zYV/U2s06eyDUzjeEIEDXbqK9iC/YDlpbwvIn
M/nWCsFawfia3ky2mfuHIYmP0ngB1Ztj/JiwljQ0cTgO/r5CXHfPb8aNoNqw2AIFyM5Ep0nQKs5N
xA8qyXfDsTnSrHs0VugOHUg0SvgvgWUMgpPqfATOiYFIrj24h7o1dQci0djC/zMQ2eWUP07I213R
EEn3x9mFSL1D2xuzm94cQMd2w74G9HKHySDFgOOG2Oa4oQ7pDZWFGkbF6smBJsXkW5A0KhvD/FbP
wbUGTkmZFmhcl3sU7t5YyLqUDKeq1uM0g1KWpF9GAdwJv+jzS3bQUg2Ut7TOey7DmrW3OnScErX2
3cI66PtV0jv7X08OjTcl9VoJ1Y1YfZ791nXLFbcRcv3qiFwK8Ofk3udbzO4b6Q8g5Yzraw90RPrt
VWZqh74xAXhG2XMjvNxLFHT5+u5AIYMAJmG4+pjNPJ5g409iAGwDR2gGxFF2Gt3OyEfOPC7dH5zX
AJFSQ2R3LiCLgDirwZvYXxRvPolzy2UVShNZQ6kXJrn8Fp267W4OrhtujS4B62CEcPb8xbDTuU5I
dmo7I4evjoGVm8reFdrqEg62O2mw7ZVjflG7HnbMGVE8z3Qu5ZlPNKWUG8vIc3rIMkvtUSny6r6H
0wHLaDdrxJk7PwCuyRX+vvI/IWFPQHxaF5c+zOzHwY1mCJ8HjEgVVbT27LnU7O0pz8sp06VMw8S1
g2x6vxqAjgUojingYRm/1R7aHmEBck6eJj9qEsEQ9mV5otliMPq13kxKPnE2J4Z/RyFm6hSPKson
vlHuxncrFd0vAyNe74BkdEi2u45V6g1jC1OSp83ZmSzm7HE52P5ZIsC6Z5/7lAojOMgggnfE2KAU
lBt2oF/FdLexiSahkK/FptB3gUh4Cia4aCGyn9x+M+K6Q47ppOlqsj+Eb0L4pNliYrvYWLpUZ309
FBtUkaiekZwlliSFk5Ux/Z7PaH7iNCRcn4FrhF3sk2NmHWoU5FjDlU310XfV5Cmmqf9Dq7oiFGbI
+AAlh5M47pFFEGZDSX0cbFrsyAmVSV+xqw6pc7qC/M3veeRKQe1XMyVwg+dHqx7iIP6024oV7n4d
JmXv9O2W/8gAN0pm+vHIdKDQG/B442SgIu7dEkBUdXI0VSdUhIgxO/1LjaEPORr974bNfgfXrhZN
vG9Y2Mjm8gNgnPCyxRTSCjDb96Y5WOe0YZ4c4qNg/iuvBxmW/myT7gXaq5gc2bAugZEkrguMq7uv
4NPdqdkE4YF6MUq+vIGEyZbLhhyVs4g9xV4yXgs4T6jXwSE9Aiv2fNftojM+oWLeh8s0bkBz6XAz
/yJxEDEaNXAp2sw90m5VKiTa2VbCurMut13q4KyM9/cwXU4yJQKelhwU1hC6DTUwxJp7ifmlOlNC
fDiaBotiCs64eGlQeSySanrPhhYmg7VPX+S25EQnehoes3yuzrCxpabEmweG3nJpEzvINdeOdIWa
kNpjU1c+V2kgtIUBcStEMB8JufnUyiX3NLP/opjcBNwlOjrnzRjKQWAHtO+ZY5BO0vDDfO2oq5ta
iUo5tJhb6UIdyILNc8cOWViAJ+levqzNVXQ/eMEul1E4BbRxcXE0v+w8GRCoxhF1VkFX9pwlB697
1lsdt36nWIGiD1VQxZoeNFZbkRbarx9AAIa91V4+zc9PGIZIgYahjeXt2VrVvj6zeHzebqXdnBiT
YnS33RCqBCHTPMMNImEeRcWTv8iK2ntW36wl0yF68UrlT1L0NgIh2wOtfVR+DmzgEOFLBZQ6Nkrl
mfWmCBA7se1Qa+VL4uyIjxCBdqxu/q7bPLdfct4x0pFVsPzH3zAcngwh1QiJfJWZFFZwUy3xsBqy
PSeCj2lU6BRd6+EiNqUd4PU9u9fbIHnLdDSqdPP6mLOllkLcU/0HzbVnj1+WrUl3nppVKogmlFUp
+PG3upmFFNifcJIx9exW0jr2pgdwAQ8cNER0Gjb0zZzHaqS5G6R8Yh3/XKEV67j9wyIGCaPSKtHl
FpMv2c89JDVGZHjYCDz038b+PSuCyTLDea/EjREfxOhJIhmMlHEwwjMtUw9Sx0MVTy/Bg6l4t+t5
MXwUdPOd6F/hH2LNAVAOemu4DkcOaS1BuediiyDIok/cMXCHzbWHAPHe8Ms52AtYFDxzUnbBmiYK
OgvNnZMiP6zxnKxOLLDcnS6vgUbSoXsY1n1+N7eDJA3LYA6TainvA3QFXZCBfuKrgiXeMxcnn/VP
hO9/kE/cmVIy3i/zKXK/4sBOpbD7eU/rUVZ8/Y0DZZsfZtWYa1HqzSvGXanQX/0pwW/hXd/IRXi/
ebDJylOneFTAZPvxhdC9Rx6hpCLOa6IdAAqyww20fOGTvxr+xRUUSclYH1X01GRH7Lgpd9XtqpOn
wo6NAuJISd/SM92I4VZBgFW4ajDn+PSNwbaRX9LK5j4/kPukN52i/SfIngw45LmNygDiFRIJ44fu
JIaMkfN/go6Lvl7YSzSXIQji2J3UXJAmUBGFcFa4Dg7B68zm1DndC3szJX7C5alLSc5vPR8Aixdt
0W+oLhu5aQXLxGIVK1lQ8tLOEpO63uD6/XxrutQluzLK8gkhzDbIoDX97KgizJPHJAeocCHBXlYl
LKHUYYAwli/iLF/W/LTGu/y0abGYwekAH/KVfm+pNq/OE9N6p0fk4SSe58AL5Rn7wqyAed1PVjQ2
gH05JYxw0TGzJ41shdFwHzQ6p/Hliv2cEsl1pyD4N8P8hf7i31vqDh3pwMf1IVINtWdONhBdFy0B
04b1u1bIq9GfoneC+opnioY7Z7FRRMGhGshIX1FbMAQPT8J+HRnyl5hM5kNNqhhf3pkZChlr6GV2
G5m03JfuKQaIpWely0hNNyVc9Rhm0hbsfi7tcBXX7LTIS94lpUFGR0IdEpbDFKnb28/dh4nIUyHO
iJ3upKLOtGqOWK0DfwB9tL2EREdmvSDXOG7M6eEdTHTQDe90xO/sO69rCvK0YKDxBc4Qv4Arjk4Z
7ZwquXm/luCOiDvC9VR7XkDEZk/BL/SS1MVnVZzG5b/BNZO8KIT+nRxQMzZHemDXbCaoIAvgjTEP
U4CoYZYItG+LeU+jtse2I+4PcZXpMWi7qj3Am1mAAvl69m9vKwFrIpWXSMQrwCeyJXolrAmnz+DT
7tmoqwyHQj9oZ5Q3TBarhWRRGdOoO/q70oL0Dv25a+DVrW2CXzNosOagEasKcbFfAPTScI+ouRTA
4ibwGLW7iErSZC8VajACszgmlqSxAxXtImhfMTM8osKKGWc9ZtQm7Bc8RbKs8Ltbu/WhdTd2z19G
50CtVfM7y7ZN5UiczxAb7nzgYw9hnQuGEXL8GuCMEWt1fYCeOPAdtCMXoQAN3XkkeuNBdC3MTxIC
ntlUECieIvajwBWN8q2zKGItwlrOkkLXUue41tdhEdfQm+E8Fi3G5yCPbYRKXGU8wlvYFzz2jUCl
PJa0Gx37kmDggT2dqwCW1v0In1K6i4QhF65V+txo0xH6YvAxvJSw0ZtDbYbjwCE9FEK+Ew/Rqbw/
ahAxqhK4wE21nv4L/u2G+xFWFH7jdeFHjggKa5ktG0cyepcRjTEq/0CfhIn13vcfUvObMdVjYpjy
TBC5wFhYrMuLoZs6xqFoKrwYdTR2ZaGfNKGhRX88lPNhLzLlj/Qkx7Tal1PA/ZP/vQYGmJtDdZl9
AWJUFiJGqsNJGZIiDYcNtHOe3q+Zcm0BE68O2ieKX2egoskZerliL69Dmm8BIAcwOyqkgl9WGtsQ
yzlrt7e/fF/qmzi6gS9qBV9rbAvrivJnyT9Ps7obd92xk6DkHWigGT2GuzPIQAjRIHbCyhNoS/wP
dZttgQ3JRh4L+Fy3Bm3MiWfecqijhUFTc0uGJSGLCD2gR6XNofr87ydVc+C8bid3zCLU4l7EBPPw
8dYuSdEfYEKdtBRCHQforDOtnS6TMfNPEGyvB49zVH5DVvBx/93hWIQmVU5SRTnoEAsSszfoCYwK
p20ZYY2fH9HRg3CG/hY0jdw7ioL42xQVzmsPVoGfQzhUZ8wWVoWWF77Vo/IndtpTDCrmWmZifPeY
DuLx03d6evVg9MoLo+YBcUVBtiAu5zB0Z2mNi6GhJ5lUt/h3xzs46Brx4Olu0u1hQkj0KbpIGH30
HkeEYPBl+UkCevtG6R3WGRKO91lcNGVdmB5stx3R0JnjZvOFvKXecOyRQlBb7qYY1sgCHq9fY3Ej
6B0GtD7rnH+ThZ3r/5KnAA8Q2H20BEdktNtEdjeOEL05+WNYUFQB8Alpg6NsojfHqTRPYWnm4pBX
7tRRO7J7FIYM0QWQGT23+V1G0HQVTE2/h8Ug+mmiPrU2731JPnzseTS+O9LpBTQzLNE1He4i+YV5
h6r0JJIFehu/59oiycFXKaIvwFNNpytN+mbKTOf0gg/RbQY2aCx6JoHRoOi4G5LXA6xZxxXbvnQi
TOnA988+N+CKOaGMfYr14yLJLQoaSXLut8Iz2BKugnKEPZfEfNWBQ7d+bwPaL12cqnhg7zcqXwWb
68Y/bQnQNms6oMVoL/61r6WXu6fJGlRjDKlAxGNE0oCeykpZq3Y//vYQYLHoi+kqVZeKozmtOkH5
dYrVSEXHsMB9rKkU4hXs0EVfIirzToO42iMJY/GKminhMaTJ6QnT70HxA1nm4hyZcSAvtkPO+85h
qsxnDGTmasFsM7AvFO6imGFQ4/C2Tl6BNXnqCu6qW1CJ9zk2cc5wo/gQ11yqZbU29X9fcaNzZFIN
k1EhbvAPb/VF///KjiJoXQcu1pUdR7Pa+yCWOvs2BbGwafjqGnFxUdq+lB9ZIBkr/hzd4/EJJ5F/
Np/DjElo/bs7/iPSpMfQT/wM1uqWuqphgLTjN4f0RCqfeTxEl3ztUMsJ4tuswxZfOTibkIwDulJ5
/C7YdHyikfFispLVBn6pLZTuS1MGvKsgCy7ClaQPJLl8F3a60FPj9EwE1xGhKq6PN+Q6FadBLiWs
NQuLtMkTvgIHgBmP77Pp4z69B1GuXoEbFNMdgh7ecTstNnCPlSfDH998E8+NH3SwMoqoTuRXtzdN
Sjbg4citI/niQyPlOrYm3OH7IECf1/DUQ34sc3sq6a7MnxZf0zQjxSB3E3BEroltvsUf7eR3KycU
dNFxk7GYgKHPBUH08FATUqnUbUaE1xO1fbkEQj6AMng+bk1AAdWQia/5f0Px0Oo548bn1584xAbs
wKlbSXj6V3N11Ap19rrMfgyWULrYO9ih2aLdAgELN38S3AFvzY6RfUklr+LV4pLo/4M2LY7GjZex
msdnd//+bhgvjK085BJqlBKdfeFkKlqwdR1smyeR/k4xNMbuwbbAHjCAE5KhBkizlp2OEqGV0nKG
5zAnDlNP1vZiScisUsISWKVErpFt2eUBFPxqfjEiOwlSsj+5hpTGl1GgNCVfGMwD/TnSl2xVvHv4
PguluId6nnCnP21DEv3YsXVX+qTPm5uRLrHhAKF9G3iKJjMeghdWVxACEF2UTK3Cx9a+U4c6p26a
5J8+lKwP/v3cSwdw7sbtCduLZ+CeYtgkCAK0uTkebyYYjfA+pWsaAlJGtwKhy/Tx/Q7yK1jsu9gf
jvTS3CpCoV6XFZW9ge/Rbf5vWXQOlZ6QQh0lAXR++jsjPITrLcv4zYzxMdvc6NPUoEyocUfSYrwL
QdWuYYeBrULpNQSmaPJPxcg6QHc4GGJydI7KnFg9i1FW9e3pUcT+E5AmVvrM1PM6HIaoqcrToy+o
gDZ3BxJB4acNxHcPO7ypj/61zWiR0PELbinn38C0Ie2CIw/fMHghlpvbS48HYzUXrxTWfJbrKrax
J4bQU6U1If0C3xR0VuRgRY07oEy7dbIYRelUCcoXY6wnXd1PjEkTLlB9ODlDFBs0v39POKY1ugr5
6gaLuXemmxH+dJ/Ul3Y3RU/OHl4Ku4vimast7qqCZYBce83UiWawfIwOhyuGwN4nZavfGt8Jbaty
+36ivwhXjhVSKqxjuRm9yhcAr5GZ2siGXguLRb2Sh5+KiYefuOwivuC5cLpCvlqEidYSbSz407KW
0SHIVOHj000i+hIBd+uuCZL0GcStbUWmSafc2C6jUhmphQLZTmTWT/uv87HHSvsZHOo3ogynJ9lw
++vh210QhdLKK0AqCcYuwoLjKVjupeLh2B0hIy34yI+YflSCUg+1h5cGbm39nPWDF0fjiKiPIkh1
9Cp+9MO9DyOqft3akhuFjCgj40zijz2hSOufr1Q2sCHu1qLv7kuAw2YV/vP5BkqfG59HiK2LoX3q
4VFy2VYONHsJw8pG2HsMCJ5Pe2p7iTeYdAIG2aa7VooxCl4AQtg8Rv4crtygBeG/jDoDOd1gFp0b
VHakISp4uqltJj58IaPstWXYBuzn7f4YhIVNKmybK+fNTQHlQbXWpfcvqcR3ZYpyY0TT9w7XtLc3
4XhQ1IwIJLMpKryo+efsKLSDMIlS+/0tr0YmSSirCyzyZAM+ya+Jp5p60XptI3ykdt5qn4ygYQm0
gKGJG6DnkJGazcVr16fD7oBDUMAMFgUHGtwc85LGVQEc5UwmXcDtpEtaOPZOEV0gHm/hcxGaBIOF
QM321Ox6w+Jb0KwOzj1oUGMZ2escfNKnHLu5TAGpztviW66ck3gcb8zlrJQYX4pje/8yfHyG7Kqw
dEDtxR7mlJRogiIK9rg8j0iFGEctyI8oj4XcL4HqLcGNainvBKsVe8knAvGHaOABCuhf+EeStCpy
TyFGTssKJgsYB1cut54dDlm9Zs55FTo4jK0SFl6I1inH0aYOVSVGTYCWRrocbuqCmcwHPHGM/pyS
hOCdAS3TZNVx6nkiurEPidarBtTFZjlMOQiyH/XJtAv2r8lMwgrl3Ax8CLQ6vTPoE+r/a13VVIuS
IgN+BAYi23BdiCK2X/FhTevsyG4Vk+Xne+8wJMVJqBD3UOY/A7tt6rTo47o9IPJESCeUg0mpveJ+
cFAfMem8bjidVnwdhEM7F+bLrXlf+qcGyjmW3b5oeThvmD7hbEpQUkiCaXQETIyRGsNfNlrFGFOv
7vnF1ryWWzPh5Y3BlJxjv8kjQlcDP6Y2vw31XnAM4VVGSfRj7A7/pi9o1CYpmDxqIKznSt+ViLeH
7cxRrabdIK2Z/CQ//YhXS0HxXqVaO6H0elSsUA2Ok4lYVIdcytg5MQhln+sj14a1p+xGnK1v7x5J
nNAyTLfPWe2aO4cSaVrOFv+O0pcf/QJLDUWNKrIiIhoKZZzqApPlNBIvoP7Erx0mLYOd0Zuk3vrB
xME3GoIsDfHjepLqSkx0D5nwqbOrmmC7AzMi3QJlxJ0xaTvpmOrV7foudhwiRPqSMClCIkUKwRCM
YOrB4QOJOfnl26oLDmWYFtTzFSJJAAbQkvXnUcjgh3tuisMs2H01uW1AOvaLoaEpwZo0U5lpjDFK
yBtmnXqzoZOlMRYa48lMf2zMGzrenm6j17BHsoyc55hqQdFFZ9OXQvF9VWxHdXMWxW57Fz1biv2E
qch9iyEVToVba1GAtOjXIJvtdTcR+lTToK4bc9QfO+t6HMgqpRUqoevWmeuCGdtVwbhzaYMGVZWt
gmBuftpj+7eMoSHUeE6MoAFtLyJIjF1fUCxMWnWvp0miaxM+EAUAO4P3GhiN0iagypEIyol4HxyG
+ilDgZK1kqywfPdSgZUBCmS4ryO2t2JgMqWwvt1zoWNzVVf/ZjI+e0jwAXuOu3kcemMUxsT376oC
6Ig2u3+kax3lJo/wr+7G6pOtWdKzIyZIwszzkssrNBGBawIvp2/BUtQuj3uO8ivpA5YKoZVfQGjT
pHbpNQMeUpO+fOpQhTnHRffpgbTJ6c9Qvm3IdYzyWW/vit+uF0fntBc4BCZn+4kA9jT6hwt+c4TY
7dRKrEb74Uh9e1NWmo8tzjwP5WjHVZyyas2CfmCWjWJO099haOzEvrIDq7tVTZ36PMvz7jikUQH3
yKb8qY4iILjNHEl1ISrXsu/x8SJbdJVmv5yvT4RxWASvU2NcjLFd6Tm3Dx3fMLQZT+rjtq04UDfD
Dbs5dJnvKsgOgBbS26X5mez2wQZugsbIVqG9i7LXJ2yQGc4r9l4JRQnXUsNl83IuP8MDpmodkD5t
5KTVYQ4dS9Wn7RNk695AZpHFh8aavZgI5ei0jxgOuh/3cLlHIrb08e+IiwmD6CyEFvdiwEWeD4Lv
h3WdfaCV4HoS/gKKzOesjEF3iqAKQzqtm6qBq8IBxMjtbAfmRSvMszBqobC2mnduMiOaunbIfhB/
+0EGNjkvEGkKRWvlDwBNRa6rXlYV3rWJnlvNwqx/zzmgNzCLaaF5nhSPUIr2WUAv3ZTQ2+1Ewhyo
6feK2oQ8Y+LIj+cgO1dLhp9JRPztPNYOAzu8AfGWqQ82mJXmvpzxMgLGfigud+DH5JEiswbHylqW
l2IWZHTvZd0gIzI6zUbBhwEILLZSPQKZ+G78dzfGd4dqVJGkiGKOF97qt3KuLFiGRXm0VyUGVVxG
xkCiiZ0VfR7g3AU8RV5zaIfAvdc8YwCwBdI62MJO6D4NhCS1Ny967JJZRLgl3lXdSsVWiSRYfODA
LS3cab2lzKhKuUlUsgSAbJr72DGOw+C9n6OEolOh66w2oKY9ERDm0wmoBA+ed1qH9HDVoULlxwb1
vT/+AjisLx2cmt0PInxhcQey1GjdgIRWzZqCZFxpGn4cBPuJiQH3ZRp5tLPUhDjZMkTmFV14Xund
vw10B+/p25yn8nfku6Z7P7vQZVrqE3AEkxGVgo9j/TZLcN72l2MY0dw6IbCda6Rq+QHc/1O5KCpF
TM2xH+Yy/u4PWKtjREA/HP2y/WYW6nyB1+FpCCday55tn25AeIt3P5x9myYExEQVm7jeVeBcXxme
Lgi8DS/fOZJfpc5jc3GGW3PEQwfsDPTeMhLL74XyH9jyAygdi6KpVChwEU5gElKcv0HpL2wN0IjH
Gmwyx09DSVBMOwiJAuIiGVEesdn0eV43Vu53gxGKDrotXHSKGOEsFEQ25g6xKxpNCTmS9k11p8v0
XD2LOqYtoDMhUempmFjDGl+H240EApjm3g8aGkoXnv2pCjZ4GFw6aFs6UN8sDcvPkb0dmQPXmwLs
Xz5Km4idNABnd0UV2DUNewy1D2IFq9mPAGpbOWgQRAHFA1mjMX3FGRfeIjso5c4hlRlLiOedr0ET
auVqa11IS2y491pe9XOM29beA59xivuCaEVYBjkW429XHR4EJiqDQsh7qnCAuY4Tt6kuWD5z4rI2
AriaAWbPlN0gy8ath0zkQUL6FNl2OoMjzCubwJdVWdPCSUvuNQyMGf6nUYBy2FwKJa53e+Qm/pgc
Pd35TO9kk7ZCM+kuDEGdGp3E146Mqk54+yDdwy6x+C1rXWqN3IghFhEAKp/DEEbJOG3MMt5YEN/d
FQMOWcX4MM08389bgr0o2KR5asXY29evcC2AjYCE0c+1V1GnCcnxPzE/9T/P9JRv7mz/AY5J1um3
qQLHaJ9WSFAjfOiYPUSWg30+9r8inYGhGnHI9QmOSJYf8vuR+TzUbZf1t6fj9ydT+1zqhwHR89B4
oqYtEGJ+s8GHN4OBHpZJrL6LQBnepfpf7W9no/M4aM6DpNfcnm++OIMdFZ/e5MjgSIzbWBp3KouX
s1VE99B43yjy3uom1iU+Swie77hXdTLfTvuUu53DSz76roo2vPhTKkSocYuCfFsHMMm30OjIHabj
3cp3RdMIlx4JCtp+yRP0LbflDLabHNjUWlopqz1QRd39mNuLg4Iidm/1BIXD687c8JP5yty9biJD
1BzKgSBnf5JNL55kMX4WTO1pZ2v4TJGpLwtKROEz7gTdW4JVsQ6ZdpSNaW1ZbnnX2cXPGmQIQT4O
4OtVYzIoHq7y8R3cEYu0VU3zQzikpIXB15aRAKHkOt6N0/PeLTB2qI22UcRW1El1YF/zqJr5eEwH
NFHwvmLQTt/v2+7NuAMsU4Wgn0KGm0CPx1x1nbvCOESaCeCOGJ+k1NG4LwD8atMI+YCxe8U3ChZk
/gBWfYZzEgslF65a3vaDXXcojuiOyvVSxZPrgV66ftzr7llhrXzkEsSn4I2glKZu8SwzqjxKOZtz
G2Mr8e+5hw75F/N9YYVFgym0gnlhFmiQclhL2xegFodZkKB+frGeEaSHP5J9RTzFPn7hxMGcKWCv
Na2uJnWUEPWmwIRsrj6jEfcza/QAGhtXaUQIANrgKuVylKcgxzHQTEI8eiMCDAH3MG28B50szmlL
AJPJTcSv24c9lH+1eYIWXsRJJ9lMTvaxd7lOXLp6T0smh/Iy84QeRreH90pMSqz4RS5BEMkj+5RD
voX6tQYTZOo7Fc8Eo1a6wj/eGN6PHpN8OPPasrlmCrvX/KeQGIIlgZZysUPXYdrim4/qeLW22wae
+jNcIGhJKF1kCTRgdHjHaFNMh7d25F1OKhU4psmOZE1ZjLmM3u3GrFG4lG8paR1yI+8UrlI8ERXn
6BM30fNU3AD8JNgahUaT3zqW0l34AeBsQ0y4cdgKt4FO9A7lluBmD1zz/b/SxVOUiLE4hkXnXstT
4nSQfFXHCo8AimDUe7ZW3kbdxUX0F7u2PWs4p+Sj99d61YATlty5eFRzOMILCm4JgBe8Jdov/xyV
r14+j1Vo5SLia5ylDwYTFH+/w5Up4l3gx7ZIbn0ICJFJoqJEszNsZpJdRh9qAPNuz4fHB8hoibKO
Rk5zbRqEy/vK0vfP66Ljp5QoMHoFS+U7wu3biYOhg3zlNeJSrtKszeYKoJ4QHDnb6c4lp48UxYw6
1T4w0wHrYqnjECnv2kbH4+XuxEVPfHwBtG6YDEaL6XrEAUe/0LOUn6oiclfDR3yb2eh1ciBiI0XB
XFcqnxsHB1d4/PUupf4oFOwO05gJwNoKNK6bYWIZ3M0xPYD7mlHr9BLK+7jxzmqRiws3O9KGt6E1
C+airiaV5+M4VJNur5kMmRPTgNEpHOXPpIvZMG1MBK2NUxHwg9lzYU70WaZV3nDd+n1QPaX9e/JR
4j8/l19dL+D9yvX4YrSpftnUP1bTbrR1l4m1TdXV7k6BuKV8jz2qxyF6DNV7s4I+5P90gskb6D6f
1/v5zYl2HfexnipCZVoPAp5+uitbPauNSm/lUvY4h4LGVYc1F0+VQvzELFeZdbb9KG+XbbwzRHfi
Pm4uYNOEx/pCE1Pd2tIOCO4MUeFI+Men8KzsEgaCLczM7ttp2BLzG/HXVOK0Ba4BryQQRK1zyIen
/Ur3BsWMHwwsiqyP5UmDykVg/aoKTgIrckArFiFwGfXE8KCGdI1n7PdBe7uvWTWkmbleifkx3YH9
vg3mAN4yFwqfa6xboXmmUvwDnpYjzJKnEs7dezOBDyUjAno9pJKyYVvoy3MHYMMa1cRroPreGeK6
qm7zPZLX74KuiSyrBLB0LRiKTJLtQuYGKStaQIzzdwujtxrIHnKKNCjjddwSk3XF5UVkYm5scT1I
4+b0i14KYZIDX9cKhmMB2hLrXWptjO2td6d9538P8D4Q0y0lvQueb2mb0vKvi5SrDdQLtg2Q6qUK
GkYZIB0l0n6hz+Bv75cz5dQniBdE5QojZ7eyFYZFi8aKB2mS9P1UbazPDFJZ1i1WlOhmncLNHdh2
oHRPiulxDhEELk1UtV4+UPP0r9poGULZMXOpDIlyiAsaFLrn9L/pPAsCEo3kqAfu4uU/yzXfCixV
7qTjlyD8vvupAAPQYr5X2SC+G02VLccym9ofYlu6IEzLJU+h+4NWOIkhVzmSrHoicUvxOa0DbJgM
MJTJNtwCe2Apy21c+36enFW+2ajrWkiqtTx1cOmaw6sbi0TcTG+8fyq7yrVbWyiMWWDMnctSORca
H9G8On283AV3lmvt3k9RuBd3FrSTOR283OVup3Bzi+yicD1gics9ExqS7rz8a3bxpUYnS3ZDtVLd
GbM8vRqM9hxbfuZ+5p7VzpmbSqWgcsv8ikZYAH4UgsxvYWXo2pOU24GbmBkYxQR57Dr/PfZ11Rp6
6dQCx51sIzvoOrHxVahPUa6m2hkn7igcKPCfTH86EABt/5taN1fG7B7R6c0BDWgvnYYgVwt1qzhO
9yg5QpYHkCaSTFZORI3zHFo/P/oMvGaKYoY5//s+k6IlVkeRacm2LPjhjRRPaKn106sPv7PzGudd
SnjP/wjOtthNiRQE7Xch84RpDQOGmPIqvELs0hT7P/1IJFBSi8hGxpjzcdvP/YjvFnvmYajk1ou9
wpxJ+MbUkQXrzU/b6z9pC3FTeAtpap0teNmg6/A9vBxGHTZ12+tvu6gL1VOPGENRpNo/4bNTtP9F
u+zxR8y4lq8ORyRgtRBgynDZmObgQbb65yjjHtFKKK0rgag1doUMD50EG/ysywP1ic5bJoKy1e17
0v/Y8Ez0H3jSnT2QKJraUVKNiZ9HG25+qvIzuRX7NcmN8hOEj0sQ1b3mcUeKsmDM7BxY0R/TXb8n
KaAQWrzoXrOD8kvSgTAJUCfLOtv9bz5Di2c/NUtssnIZAH5o6QL/Agt8TqGZiyN0EYNssUQngYOm
jCVmXFLN5Xr07HYcy/WVN8elcZ7nzxEL1Ff82BNuKl18dkFOHEtpkuexoA+G1Z0KT6pgW4MVq7/6
pAEI/zOUw8F4lmKnWMHjUuCIJG+wfcMOy19ojkK/0FeF9wGFVSuekL1rH0W1/AP8Fo4Orf5p9vwm
GEKDbFptoOk1EUOSIKNanunIMf5SxeNuY+Ib3rKbynLVl8J63Z1ET+iJtNP0hJq9fVfPPwfUuOiw
9P5ywgZ8dJJY80PN6fCo0xFBpmBqsMcq/umDt7x31tvx7JUuLZDlyvc1YyXaoEm+SBXZMn1eqF7T
pIgV4fvXRxXN1JgFdoJGx+W0IUCmYbVKxF5GRgIksleO7bf1W7o4zay7vuYnukx4xcYfqCrnlN+T
+BOnE3odmbzPabTVvB1pPUgBdSPtJeDYfVaQnKKV5uL4ovU0JLTBSci8Twwq/PUbjljAlbsJ3hgD
HP4MQThtJb2qeMbKTRzEZxjBcEM6sKa3e76TOv/OKE22TUFa0q4aEDutsPSYVl61xtrsaYU3CqEQ
I+jgjzpI++CPy8qBW22Cy9tqG17dd8r4hpsoV35uOxEkfEoSFxgREedLGNp8nVkP2JoZSnpaP1Xe
XXZkiyTeNk22Hx1W3pmZS/1UeLfw8zTo+Ug9Ng1cNCl4BQimGPD2lJiC1yBdSvnW7tBpCi7dUl95
XZvSMhU0oJB8FbhERMTwRdDZRQ7YCQ8XzBQpjoo/0p+1V7tBAATQFcEvUqSrWNXtioJeLiJRIxHm
4YkCn/UaZ0T8n4U0zZerogXf4C9MsY3VYuj5hUKC8a2vsO7Dq7y3Qd5htfnpBoguH+BlA1ATcVsF
SeYwcpg5KEakmaKDH3YOKvc/Qn0BbzJCqpGRvxg3SjY/6zhBEIKVjzbAz0GbVt4aCq+7nY0gL3B9
T1mr+siAkqmKPz1VYs8uQrPDTsRiPsxvG4U2XEcwg9BAmytZMs5tIyNbu/ctYCOewYM0GyFnI6vJ
2/iyiyoKtpQIORkFV+DIdpLubmhTY5QuvMwoZWI7S3ACSSKOvdVxsiRjSCTYPlIXoChVAzxhNtCC
dK1EQHIBejRQBA4CoLWdRr2dCJEWfyj7uZNSFYIP/kc3PzJiq4dvqXTQMBUD5bAMJUC6OwqEmezG
SjXItQyYxiMIxdBFcFkvo9BqSetVmD1lj1Nx+u390IJFDroQEcwIvmIR5Sy6SLa8G7QZHVZjinpE
6viiCQ6Ww7HIKldpMagwJ6ZmXc+k6Ux4VXyOJMB/Qm12Lq1rDr8+l6pUdRkVT+kNGsKjrcSoIQwP
q9f5zp03f29RzJPVCZyqi8DPfKrFml+atvrInkiSp2w6ej4hpHWBN8ix1bqwOegEYD/lKQgjCBPW
S2glrTN1JWFUo639cFbnIlvH3WgjucacLTlIpaqytM1iYRYv7LrTvCr182D4rbT0gtTbFnPw6Czg
foJzmHOPmXPYmKl9H0JAxCEAGvlDBkHwdj3DymIzcjJaaQdD/STs1yI4ie8zJhEZKOiRQh34Fejn
+QX01l8ucnLcu/kCnP48Hl0OMhMx6UpYgyM/NXTUC+DRbY0aLioUHEeQnYo+Euy98KWY2yl38jxy
fgPY6592G+82j2Ll0TcpkTA2k86ptz1F9mXrNcQgSpvJiV6L1bGX2L695iHGk9ls18M1OYC7jJZD
HxaMJgFb9r7CJpUHGbbnuR7qMbMQUgZkK25pA0a+jzKDdlGKWy4deyeGVzX1WIMPDrDuuj27E1N7
4F0z2kGoerjw27KsNjDm8dRZTQw5LBdkaeR4Mf1IR18k3Mvrdt3zMo+KQfCKV0b8+m6OejoGmvEU
gpKCfY01RSsMLSTa+80V17Yirg5FZdaAPrzxGZsIkKQRc0bnkV8D7wc4mSDPlMXJWn0hoHmhHu5J
tlcfSQk3Nb+IREHCD1GrIOuBeIzjcdq4+8d3+r3Jh0WM6RrxWNa3j9Tr9ZSRFxyLjpGj6QKQZLz1
zPV3xrBPvN38kKXr+y/pWyq+y7v0WOlrLhIWS+c+ZRfvFALxOHKAYP3nStzpu/4k5TA1gTEUZEOH
cuN4bXUkwntHYwRt68lpTyOG+tiIHlf6zAGko218887ocbdCBIIodk7LRULdKzX3GrXI/nEAE8RX
nhp0uPg1k3molrBATN0gV1CtnmOAVgy3zFE/R8lTYu834prZQYul3PfJQqxZPzyMKGEFgC8HezGr
G2E1Xz+ExVkk0QOpEwB1A9x+4XiyyJbHrZGe5w68Dpma0wgsMekD0z6FQogK4w2VNtnj9pi29Dfz
5XxxVa+FL52uu+cvPEj2Zgk/pp6KO1I1m5JP60bozc55ydSlqagEZLZq2qHI0hw2/4i331JCPbIp
AqAjgxGpz8sdAkSlkOEnhI8dLzeaZzFl22docdzCnk8AEi+5U2zll8ENp36JFD7yHkQUkbDHGMqf
Mhg3srMpXVuZNhCwwoE+LW/Mh7WG2YCEgsxQvTOkWbHukjAXwQbhZjXEZtnCQdRebCHF6bpTbB81
WIvt77L7VRp4caHN+GJSuFQMlUrK8aYvpN4R/B8EWtMFevaKA1gzREpyXvnfQtOr19w0LSidOPdw
/1bCkHBIOnKjolL7iPQRv3cFIDLIY3mes5ziyeMymtd4RMoDaH1ReJdnPNhL5oQ4LwXzRc/ZCpeF
Pm4mrL+NSR+J9jXwQHmh3jOu6dl+RViu/w12Bs6kUEGzOr4FbbsTIkQ8rpmfYurRVn2mzR6COQi/
qAu7OnBHcrSILCigDD/RbifPtBzG0+CVVKsk+q82iKRfB/lZgKDJUriQ0TPtHdrHDRL8XDfkTaHc
O/DYBxuJAcJ8xXrLAOlYaSqZmMJjaZudWfZy+NAgCKP1XfLMZP+VrQR12B0ZiBaW/o0EzIghDojU
xFPyZVF2CUt88+PFVXE7xEmXicd9sp9trsW/+1+/bvC+3clupGFwjGda3PjWQxdBrNCEaKCgjl1l
6iYPVJ3NzsvkI6gfkr+6LYnadYuxyw4OLT4CsSQFw/5AEuEYGK/NW3SI1+rAw5otZ2RrdgUvmJfH
KU6GcHzJtaShrYzCTcZwfHUYkXkLyHI9DnZDBWigIA8uK9g9/JZERDeg0ke/9L7rFaxcTvbDxGzi
ZZRjsOCXFw2KMl0sZ+MUleQAGu9r6vw/Xbk+bvfcdm7YowzNpnFDd5rsobqWD6hzJrFmYlXK5ME4
cruPwYXXqlmE04rX7W4L2CKAOaxqHo1eRXHnpc+6xNApSVpG+5a5XvUuMJl8wwc7PnSfCSC7gkiF
LtVUTp7O5fQFDxuwk64lx2+yNRIJLuGkiCz7+NgQY7WBzWxkcLlIoTokjf/iaDTUFQE1gCqsa61d
lt7qLcDHfQYY3Z+uivOJLky3nX4My8KlzMnDmUYOI1Qe9d4UMWZ8yuqM3kYC6gb0urC/RGGQa52f
7k71UWSV84pdAVyPYJO+pc8PUKm8l9m0SxEPgCcUvFSsEs/aDrZolD2Q1Z84LUNRc3R+VjB/8PCT
vdJHVezf4qt6PvrLsMzulLqt4QiZpL0NaXa/RZolqMloYQnE9wBKQsUQDy+Hk/jqLYTUkCGWjrjH
jz/HapuqwH0UHFW6FTqVsHC6hEFg0msQ1MpXbBOPROk3ZuWXdrtzE2x78XKcfmiop3GJ0Vq7iEHi
3dL4Lqx1JbaO01sVheBnbci3ytiX//FaZymyLXEuGo3pvKggVSwQSpYFcGTRirIDNATyA/l5kLC2
DzyQmeJrLQXVzsPH2ki82SYu7JCTQupu3sebHw7B5+xfEmyiwGzNhB64GEvSyn2n2ecWGyieXmDV
njylTqB5JNq0PMPcRrOMzXw+5G14Qmn49LYqjVXXmb0KO8gl4dfZmsMuFrPwekaHO0n4+rpMmd7d
0q1Ed7EI2hka2LlRkKncgM3/ItaiRpGNFDfox/TUDaEQOU9isOeP7afR+vV6Kw5JXaxKmJLnvTCL
gyuEHjaOb4BMPjikFbPBZHiDMwgdtTgsFjJAJXk0a9nLLXufDcu74Db7NqBPcI4kLzO4kuOgacSF
xlMhYSbFy5XtNkN4ruRxAL8zxXe7Tuwnx17kd3OFkJaXSYkvqrFy9KINpdNm17AP1fc7iAeazE/3
lN5Jl1+TQXQzHeOYK9ZB2V4wMzW5wZuzxSngnFYoHeryjxNBtC0HqCxaHi4fyepwnjK3LamWL+Tj
lREr2sXxpBrEluiN5rZjBGJEZ0NXQcUvIvBcaUU3XIWG54Qy+sITMMZ3C+NlNdqI4koT3W759LuM
fU95tggKet88yNhBaNI/gt3qFxjCOyvCLBq9X7FG/T8lhO7SP3y7AXvVXlPJczluAAr4A33bJbRt
oK04XY84fAt7jws0fFXvGPdPLhrwxZMtivC2XEBj+f27SbyaSQmyeWV/8dIdUXhSTSC3qXzOmBGn
ob+LxDSkJXn+G+yGfpHxiFuS3RZySZbtY9LIq83Ygh3Hkb/fARfzf+A/T0EkDr3smHqEMfUSPfO4
c8TPMObn6wezkw7RIL8+p5DFh0awvQeL2urxev0plQpiOLdDOUZSqs/QE8hy0d7X+Fmyk4AHhL3c
oJTg59x3rwsZEdobCwE6AFtDHhEHQ2OfOKeZ1g+dJ5H3qYNG/bf4uH/nH4UlWrn106VAiWmey5Zj
M7tva3U68ZA8A2ztHjyNPGIZA/kvYOtBfr3KgqGPvkwVqeyVHRIZuFBFxwwyZ4vr43nqZ1wsIQgO
EZpfhTrFTwAWv0i2w4uygToD0cJZlF63OXJYs1gM9quYKbwNPkkVFUm06oCq/HO7KiEIdgafJHUR
HY4tAh9P4Tsg5oevGCkYlTrq45dXfqZueSsPGZrpyCcVnIr5Q8SRNJ4gmncFQ8qJ9P1XBSX/ObOv
litHnKjjmpIGvPxRXfxA9x+4X47jU2Sp1O8qrNmV7C1gPZ6BMhy8ZEPBhbUOd+InHz1yCQTfq9oz
T9kYT0no+VRXcEV/ZpNDAbbr6RTGCjmPHagtJdADYp5cWzPVE4S5SAI3gCcrijwlGTiXzzB7wBtQ
3XyRW4X0wpyfNJaLVDM06TT4zzmkpBkZg9Z+jZeGPagLefczUAVaQi1QL31TL4FgCou+7BIUvVzC
08LcrhHxbPujUU5RVT/EljrTXwPIVYQegNqAA19zRanumJ+etY/AR0/oLrX+fCQrqiZzD31xwrd7
PuU2hSa2hZ5zOyl7oOUC45T0UXMQEsRnvMix0RG605maV+o++b04t3j+lylRYexJAn2TOIClbs9y
wFFFY2cxpIZRYLpmtiK9nsjTU9tM3/rBn/qdcPfmLWPlKZEW+BcPKqrg+K0oMTzJr6ztKJ4aYPMW
WalouFx5vUYkrbTPgt6ctwn7TwvvBH2vf0CTNbIfkbaQwojGF/CuMmMcl9wyQFvHhUyCgAUHkmwe
2hRcrBaFk3NmJOpNmKvsVvf3IVa75aLsZNKz6piuwmeAZHs6Wsq2YAUhHQzM5Djlo6qq+KIlT67s
olEr+xh8aYOgFK4enHKlFpA0bgOWrU6Wc1WEMDkyyQEcTtQ3zAEbApgIQOoW1a8/DxQ3ntBZVWc/
kQDywv3+tMbX/n8msF9/3ZursxmZELWb/FrdjeIEdhFdQNJ4ngBDw0Pgd6dbz2hAYY9WTbgKxNCG
RRo2Fl9zjSQRxRhG36DkKTvv5HzJa4nUAkYA+Hv0+esMUM1ACqw56iAMdPBVI/xp5QDl9hQk65Ut
zH1a0yZij+9ekHrrQ1bv36MzvloT4p1LN3CiUkBz/A3q1mRokg43iA4OoizeHXSKrFb5m9O+gtM1
r8J9/whjp+R/EUnP1bcr++rLgZ1Q28yb1/r5RkdTpP3+mNAXHJCovtp5DeKOpJ823uqtuwudMicU
bO+14czCsQ5k3391wT304NmPyr7Q+m192PdHa1EVTJ5QdLapVLfRaWSqT3W8Dyf6Aw+v9W7E/iFB
xJrgDvhJ+WT9oXPqcTVVWihf3TYjfRYwuH4RSBM0sszLSVWCRrAwM5Cp1Al7+2x8CRrm8DwEWE9h
6XlUGp/Srtiolr6O+Oru5Dz6qFzYvBZqHGeYISgu+Dm75J4BE2xgYhELdhr7l5KBOzZCsWLQO0Pk
RZnYIOhhMkOzq5cIEbmeypy1rlL69qCOkLw9y5w8kUNiEu1AELkJSax7edLlLdOCITnuApoiC4Vx
OZ2NpS1JBJH0Lr+ltWnkF67u1neWtUIC9meKrUcfBpYpNhbbgb68i1pAYyWjJIGsmsT3ZMiekRth
ZUKQ6TA+lcMxGXQ68wJd5eqhYao7G7igR650UMNc7/DEJAuUIRFsR8a2znPqQLJc1bmX+f4uqDvd
U100TApNLUVtd8EEXcBi55Tdx6hPMLPBzH86/hYITBezrQm+ZR9E6tSkAI1Bj7zO37LjrzsJS20M
XDT/Kwt96GDCpIqx59EAM6wu7/zOH5TBJWYe2ax8AsH2hFL4fDV4aC0HM3W9Gzx3eYxuIq+35xi2
YgmpYQwLphlvAYT9C1Q1Kop1wx6gpyX3Yxy8TRTNzEVNhYytr/RtXN8wX1k9AoFEMoe+8ltG7I9t
iG+wQUYIlHENSm55Y+tCBurbtSXxzjfAR38yQqdLtyygVoycmkKllQhvSGXj3/WEDXRaz8E1YrxP
MOP7AXCH1Sk8c8cdcFNJtdndDAjc4dE8ysuNPXVJKn+1Esy5SdL400p7men5HB2BX5+iQYIgFGuJ
yFj8OepjikLic8YZ0NHKJo8tlJT+5zqNIeh+dc7RpW7Wn832psA6yR6lTsF3lyttaT2XmF4DMt+h
quHpgV6/sas4sL6uWoD2P88/EHg9QFVGquA4cEIbXabkfUVX1L4m96JqMI6v8LnsYw4H9pCkc6VZ
kbmQh0RqBq179bjUBam9ZI+oUp6v0fKZBMzjGXXPNVFb60YgCjwMur0QxAqi5yXvFd1bQTd1VDMK
ybg2v+iy0wAjGPfGIwlIbso2dLfRcWUBqjVO29uakmBS+YGde2aTMeeylglov2Z41ZOQ8OiMgwNC
WW7DK6W8NIBwSgY/15WYhxTkwVL4L7PJaBmd5vwXDSfWZsiW2s8ej/WPhgpW6BXaAy8arlhsxqIx
zIcznWA1CxNw20ob7+v3gx3/Nr5+rYNMTDw7kyN4AzZDQjSZhUV3TvzJ/Q8lEWPblCAKWNDSIwmR
MttjNy5lxpjC3W9MLq2blchTOvbQEU5LnZtF9953jgtm9wUeTxCjBMGEiFlCOGy7RpD5wYJI4U+n
I9/O+7AenYhxkc3Sq9WErswVizXLJHhhQFmIMtsJAOD8N80YlhYknkTD9Z4MjNDSMBSubclGoEXI
dRZdgVD5Fmyv+BZS/39V70ANec860GJm3akrURsNCG3PdkDAqQ7n/72r4CVy4wW7eIV5psqgKlWy
D3De8+27rQ/cdL+8P8Lg+jLeCTUiUAPUS0kuiEdTYEO7svcIgLr+tOgLU/5GNr5kub7rMCNAyKy1
u8jsISDSph86nl7IonbRAYLtHPJnww/PAv8CcGIbJ+KujOy5wW3yqMq5QCDasVWIvsVTz28VZx5V
i8Y9Ic5cU9d94TviFuOJGjOKYcc8a2IBfTv5B4RM2nqnbLfjlE4yX3Ct+k65bqJ5NDeqBBOlmLCU
exfCvvdnI7kPf72dxDnCg9tEF/fo7aLcMzah4hBgMB9iGNA5izYBonwVkXR4txQaFbHU+N+7JlN7
i1PUY9hKWNhebGwtLQbykbjNRra7/3H94xVyKk4cIls1m591XHj55HiPZ+iKaaG2h7p2HQdYjk02
FChcgYE18VODSOWLPsT5ooTE56xdcVE6cQQqgMs+yZD+3g9x+EJn7ssNuYqaf9/zWV/GdamO00Va
JohZ9ox+iXBlsdmEeTrN4RsT6j5/hzxjYNkaCwLGLsXQkQ6QaNZ1Qdbpez9ejb8LHjIk7znLv4Dw
HIOXH3m9ZqPFE47GfT9J/MDb1Tpm5oPa9BrQaLlitqzoNoq++vr2mnLAJR99ZsCHJknMq4W9/XOc
UpYubXMwK260iDVvkYWaq/yQAXMzMfpJ/5jupSKMNdnoX1WA2IldnV91lGEpJFQSVQEG4Zcq+/NZ
G6Nho7l1x1qHRlpmkvLgB0K+SGevoxtNErbzXHqG8LEZ4bHLUF/idADQKjUay+VCjz8PVQmV1zz4
QcSFftZmtTPnVGPwky+khN/VARa4/W6fpY+DCdrZHsAuZCQOfqgRTPMCa7BHBnyCdiMXiAkYK3v6
cCp9t/R6KmS5VYpHgH5yRrNHWbcXc8KgtSiaz74XMyppS5Pggu98OZmnhCV5Puv+DvpoF76MCbD9
5YEYCzgrnSEjO/TBPEdxWTgbiO5Rdiy39BEyjlbuVfqQafftcJkPKWHbKOSnHCTwOpRR0lKCXTji
PNlzSBKlCzZlyhw0FuBWNFLSQPbIZEDWzpHWAPPS954Bp1wsE60G5r+8beVaPKQVMc5zq8YFiwXk
dpAPlWPg/Aw9FkLCoYNuipyPhqKX++W1eYlFd0WfIF+FczeYE+HxqD4gx+hQIvQIerd99Ayw1Oey
gSq6r9CudUQIv04KxRXQ3ohUnpPZYIa+/wFIRU81Lm5uuhyKrZX1U2ypSuMN210wlqeg3WtXCBBm
tBfqfKDQYiujYC4nkuLuh8zrTiD3O+3r+bNkASlIdTx4iOKOZ04/FzhPSr1ul+xVQZ5u3HbSPXdF
7wb3q07N3AT3hxjfRkBoJXef9vcohm87DQeufkBX8Iape0Hr2Dec7L1FmKUHFNrXgENjqBVqQxl+
8hkOQybTHfZHC0KvKohvhNjj2p3qi0AbUj9XN7q7rP0KbJsDk3Ho9Js+fug0ruyKcBKqSWJTZ1Kg
sx2unG/5l0VBwAZEmzB84UpK1KcJBqIJPxupRa0WhLGbSLRq/8ShynXcdLZKOJL2vFknxd1hrzNB
uZi6/QWIgNTJA1dwUi48WbGoa9MdO9L+oXCUJ2isnTjzvEPgi+BzFEHDrYj816uIQdbI7Yeq/7+y
3GKCPPFYKRzYsB4tuzYzYY2nfWWgn/S3fXPZc2GCc17kA/RAbQzt/pwA2nib8empi2kxToQSpg5c
dH1kNOTyuIA/e2uT4gB7UlZ2qxq/J5LBKoiLvRGuHEvsC5rlGIibjknr7IADst3l5IPNfaQp4W40
MNFIKg77MCaprd7x3PdjCi0ZeVkLvic6KnFcNBI5ev0SdIOBnccMy48Gz9TQYtZW5Qz+unmB2xmU
YO6Mdurxt43pQ+VIaf4HrvjJOkhQzXu6BKKEjnMwb6bc+Bxa+ZR0bs2dDH2oAJ3+Lds5gSIrpYh9
RanDkz1RX8Ry7u0MPJG0k3U86Dtoqit7deJol2qA83nDTmSa9DCXVCA9CKWGN+jZR2ymdVZLzSPd
n4dwTqhTlaMObl0Q8wgbPoExrPvs8RlqWDmOANNxKP+2ofY9fqEQxx3NQ7rq3ocYUDR0exfxlTLA
joeGSHu8A5M2DRBgRlpsPRWLaMFvDatpKj8BYkFLauYHWMwobn33xJlSWrPBDjuDxTm6L0A4HJ4J
wZtAWkbdryNQ6VAQ6Fr3Hf8G7B+04HAaOuNdly45DwoVg7ltXmt2wHIWSQv6Ft1Zv/sML8Ng4lze
ul6tYH+CCubqpY4eUPmcyzfLEbNOdYg3nDL4HZJoqKJFmk+B2UMCQM/aWxZVAMjlMk7UBeLgFXNY
jhoUkK/c1TumJGUzQ5fbuZ2zvenpwLG2EtWW/oCgFc/fqKpFcnaBPu+UVYRkJlNnmJhGEFvgo9z8
EsVbPopMk4+9L1ysQp9Sp66PLOG0njY5r9pddAPZClYAZUxrUfKQfWUsXLUTWF8yHVd/LrDqDBnK
d7JVLrW56/KQnAdi4aU20Fo2LOxlBZCZxUNGuYK6cBi8Z1Ceyr9/1D+v0/DgP4Yj0cGBSX3rnONA
dcJiGukwCQYeT4UJ13FFZyib03WEgxhEwPNTOK9LNgQ0UkEk55YvS15R+QoT/qBr1r6X8kEQgDoZ
XpFe9yWbBBmpsc6XE4g/JF2OLTbp00HAESBo4FPcwr0l2KbjyvPww1gdshuhgWgQ8aGbm6t842Z8
eHSsz6bcQ2pmbiJQ3wQwL3i5hcBV/CRIFBNGW1Z0LMkH6j4iEQlLV1KAw2dtEmekuTR+TEM25iCY
YDPyZIEv2OEeOqtdWMQtJEG1W0MP8mHxSv+6zRGJn28kOxUoeHxdRbVIaaxedLdr2LAR7oLOZhL6
bzFE+HEhnjkV4U+GpCnhhwqdvM3Y+JvCwv9UYHbYJnaTzfTYUHHOgk60bHbjVcdSLRUGTdQ0rwZy
kMuFQllsiokayZ3MdRx+Bz7SOmyWUv7Y2Jrlt2OI8/d70ifreoAwX6ECho4tp3GqI1wKl+34l4Dg
ByWnw2X5tFC87F5nKzpSxJJfWtPKvschvSBeHNhgfjuFhFQtFf+aXd1JPFz+XelDGCnd+Jeb0zKB
lvt27J26Is6T6wh+W/uTYfYCDlHeNn3Qg9VdOIDhrxwaoIt2XV/dmR9UBJ3RxLNBDoiLChcMbwpG
49TDtzovglg/l/yTUQVMRUAjB28/SDQenWA/kqpMbVA/MhVBZnKcy147Nq5gNGptReL1P1fWFU/T
2osUewa5DnpPMWVUsM+vdQgwSbXjHdmVpDmOksRoEuWnyRVhxijyPos8vpkuqjxmXOEiOPoElj2Y
qc3qXmjSw81gas0hIHP485gp/XbDJFSsbsh6PsfK1JvfPPKn0/UYcVJ1SLAhWFuB4ifZM1TE06IB
qx0p1noA6hh2qSTfgMzwaP++8lMElrrDx+ezDpvcAeUpqkcp7Lw8gttmND6nzDiXu61JgF6AuxZ3
tAdtkizsoO5tcxmYsvpzBk+SQtxLyy4zEbVdaYrsgYSI2tgvHsMs74dAC/IsF0Du16im2L4wPhTv
kwlff8SX5tzbyu6mEgLJn8Zcn4uwpIaumhlKgpP+SbvF0bvJZWTHwO1P+lC8bNVji8Bq5/Inuuk+
TLPQINvxa+4s+ttK/bQu98BssCUUfEn6W+WlLJsgYHl9JxWcwVJZ02YKrN/IZY55gHBoYAV5DlcO
qQmvcoySVFHbnqe45BImly1L+6C5J7uWWoTpTR8NbYfcRcfSMMmeaGm5HwsLtV9uT5bxMnm2UyFt
xzLbG0P7mdEKAUsd0xzvPbAhsXwwgig064sMy+BEPMaDD3tTnGhBI8RP4GfgBxtWUis7DEuW5KBo
1VUHehw9aZCIDjAe78n8h7VWxuWToDzWcF/OkTB8gWJKANwmxyIdPucVL54nWtAHe1RYKbkZssST
qMl3t2iqPFAUHQbSJOSNrx140T6zYB6+toMyi4Iq9vBOIofYwGNmukp1OO6X/SlEJDJa5XUGt3Vo
Bnh+mWQbBVutyD9IdUWo71btkCsB99G1qy43QypYeNoGHLBCRmI/5DpmxmcSESEK3nkIOC1Ad+WM
mSO/HoC8AG4PLPAaXnhgnD0Ae/GSQgA6j3cfxQeJgmqM2d3uabMOGwHNt8d6bz02fGgSYdtBKHpk
qM0ir2TD1JL65RWRLPBkWQPI1+9SeH9e4UCSmphYV7aR6Q48/kKLYPgV7BPB0jEgHc8qzx33e/Nn
EXkZbQjYxjDkjIeAOu8ZbVw1RTHNIYijxgsv6+fs8b3ol/l/jhec0riygbA6CCfM1OFuoQejc3Rm
/+0HoRlGXT6ohu/mYIq2z+ghKEmwdtnskWN82WScQqqUhVHHDcc1INCwxk7NAQNn2fehS5GOTA2K
FzHT01Z2ROafry5RkO2Egps3/QJq7SVjHO1R3b86WdEO23XNV1zRTCypfsRSfMiRdfTqQ8AxQnDx
E8iPVHk+ZMGVpKxs3Q7unepkCBngHKrn3tmQhQACeR23jHBbqFyLMm12uwd5zwjO4lDFiiuo+qOR
NPxUPp17lbAfmkdPt22Km4hLr1VyNYOUQlL63rv3uBwFddNRP/UlsYzLW4ZPoSdLmwShLbiuyE9b
jWRT6Jzw+vX17xhL+ycVpwL216Xypex4emA1lQ/4lgFp0jjLYg+YNmE5zS7s5c57ehGcwloYudKq
Mae/MKPjTbj5Dr9w5HD4TTkdHli1eohk7+LkQn2j3tGrxs/H4gYOxlxCqFbBGjbR8sV/rZhMhJ6R
sntv41K3i7zhALXn4Kgbwc4E5uwbheHrkM7bpNLaWKWs5Y3cMWDqtEd3CV/l+L3M7Yc6gPiiaCDz
n+qT9YiYrtcmlk94tMaaiclMKn9roKRs3MfGk3QQUZfUKOAgNdOQdCW/b2tAmTYnqvHXvO7ihkOE
ViZ4wq1y2Prza5D4qEju9u/iSqjSrevBMf+Ux0X7a/wXo6t2u7Lq31llwmejcBkmg7cLGdEsQCtE
j1+zrvzM6ksiYAxAGVBeQXaU5p3CT6Z1QeQDw9ixekCuPYRpCOjwx3G6IeOtF+bxMzuFrXuRwN6m
dYhb6Z+5p8W9YuEO5JuF3q8jtq0e+S+/0tT9o9VYe1vCZZeuHAI915VNStXB3+ulKlSRbG+BHis4
EB58pE6Uo29RzhuYHJJXA6N1EDvUlKOmZv3D7d9T6hpa58MBsJqVZdN3zt653MdQVNA0QeGnTAix
jMnrhyXuhTCWG3TjaW3eVIsLMTTmZUrk36jW75QfrNxDG6ROrCEGWSEGSl+KcHw5yOf8xLyCGHHT
IkVFcbhMXoYpafYQzpDIXsiQYn3UgPpwcQJFA0YuaHJLPBrAPreE5uqsMMotNIRYqYa0yi56cbG9
5hi2ge6c0v+TCX5mqZ99E6uo9w8xlSQLIGLfEve7sX5/PlQX3PyYmnqfz04tKc3Uzfn8e5paWoeA
uHv437SkAoLMGF4EfQY7Vhor14FPrukXM7TJ2sMymSRXEYhxjLWzHmbf+Splndn3lJYm1Vpq5yi5
fhM+NxskFHIcJ3DjKJ6rovcc7idhzPvWFDGfbSvPrEUzVieLJg+KGph9Lmj8eZCzUfXxeU6fiK9I
uLydUzBfHzvJm/2T6ypkVhpEZo331IYsb6CXz2yU7hV5QW5vyCgsZtAMu+iSnaaFJYI41HsmSNmj
GYzEMiELMuRFtA1ToKSZBZT9yXdyDMHxJxdKusNPJCTazd1N9iI6KBk263Y34Wsakq9mVGFYpk2C
vRr6WEXT3iD1WN2bO2wrb0inaiwnzOPRe5eqDlqIZ9M18kK0cCx2bUlPF7MosZLKCJ59rvr/vNK8
0h0xMa/a4j3ABZLjFEmP7CADmKWWNWMQVHyGQmPqEAW9Hyafk9RUtduVrzsY4vCEA0a64cBjjqsq
ZV/j1POJUxT4hblY4DqrEcyG3NUcqMAPbw1mGwTEv2b8oVL7wfgJxpBQu5yrGjvLWa+Gt7uT+E9D
WDuxQpsD9zDd3YrxVabpWH4DYx2c0oO5fs4CyLOHa8iOotkPoFTDX/VrueWBpbSJCkWZxg1TJn6d
HXYouQ2DP6WT9tH/DKD0IW4/A3KooGrnFSG2+yW6NQk1QaqWgm1DYV5h86cr8AuENn3pjowKl6jy
HlGRGmBAvcDnGO+tWdYTw5qbcHWgTFPXc+P02o2WihGQ1bq9v7PO+AMmOvrgLiUUT22u3Hdx/Nrb
m6imA6pVRAdmEBnRBsBJZv78tAL6hRJXjbOs9VG5qzaF3tEErrjyKKeeNOAgIn82Gb5wr09KeUpK
24PIJer+c23xdyAEYeJZjGb5D0twsOGRVG2P8S2W4DOXv9Di6hNSBIlNhHUPFWfYisd9yR0Hq9pt
0Xfe286+ZVHm0z/u/pHpfZBo8fGQCyZPAm10QijbnDP0bYb5TubSNbfiKWS4zyzeiMMLkcUyc39h
4iMPPR/n+DKPpX2E44EroBItmoudklxl8lq54vFZxbhs8A/Ssybhj33g0jG/GEoFTNe1zvGd94BE
mVjcXqqqI+n7DvFYk08hfbX4NOHsIemTsiSicuXkY+mqtL9H9shE1USAVsha8AoR2Ng68wk8Lotd
/eCyx+OFmw444OZJpUNSALt0Od0DvvuBM6FBlOBtnPaOmez0CO1xKyTFNFBEfjIrZzWfT3HEZ0dD
otTWacCjijzmSSygYHxq9vauWja5QAlD1U3sDCEB9j7aWXyMnvZ3SerF9XZQyHXUsfM7uccLdhSw
xSfg/KJy7uyBh6a7KvI6ptetolh70RcyfO8Ar8RRTnvqiila+57mEX/nd1cmr2tsZxtxSP70ZJhc
f0k/5SnZtWcVQRdMhPO3YJRk/SB/yrMijvuxBgOksydOG+Pf43bOp6yX+Ym/8GlQrFrJESiAZkMK
LmMTcTz477UR9rGvHB9ahzZ3c01ImdMfNL8T7evpytvNTNItjaz/PlgmdhlEetVlURzaZK1lCo/v
TmPwoSpjBU65DD04jwt3Hsufcl/T7E2kba6h2HytCAvQ3hf8QR2nwINrgzT99CmoIA8lIun8uOXo
tEmSZko9S/vyBYNxXtylpR0Joc4VRmduR1Uqc5BNVpAODzpOtYTm3i0Kn9o2uQMZyyxW0jJNtgN+
Kj/vx+aapkB80Ifgcd7wYknUNDRq5w+ZB83fjTaD3LAN/h5q6qMNQmGjQFvjAmpX76sJUCdEMde/
ZEqwjIuhlqlBrANuNmVK01Tm8Eo7eylVjh/cPUrPVNstJIKy+ADtoJiv8L2vKSxfZdRvbv1LVd+h
hPC6A1v+IlnvK5zuyoFCsLYoNdSpj4pFsFycG+k8q/eOCis0aJszjcZBtgvDHlBc5+2k4dADCS13
zsrkheYQ7xdAosThZhPO8qYEYJp9v+RSPXJKKwilKV5FrLFD37ckk2Rw+TzV84/IMMXZZOou/FSe
7CgDyathROD8Oq6bSgPcX3lKqdOXRl4kyt5pYOU3q7pyzkO+XJkB/bv3Cv7XjAPPLQekrAyXNX8v
KrYlMQYq6y4TuxZ6JaI3YMITtCN4hO1FrREvNL92EtfWUkY9+3j7kNHFeeHOrhksCMhauhZo3u9V
rqtBSoAmCBbOmTMU0JYiNjuBqoZQ6mZnCIPN7Dts9XuEQuglM4bR4/CdoeG6cAdPLOO/WZGp1mSL
39m+ufOZOYpg/xifzpS3NHS59NCzOCZb5AsoyQD2uWA36jA3FTBnZ7Q0JDsj21RarirThT0hmH4D
feU1oTmgtv09yh6e3MPXBOLTfGVUoxkOV/mycV/9uiBSVt5tRr+Nhof7Q5ZhpXHdzIZyTJ6b7bQH
6srmzJ/lEPEE03pMB6vr0Vn/vi475SeTk+Adlsj4Dd3PNYbESIqbcu6DVy9GIip8fMvdoXxA1ljv
Woa9WYcf10dHPlWMU3gc3ydBLkIzacfL2Rcf+nNFgq72OyDSRChZAkPEr8vt7s6iG5V832rlOTZ9
y5DtfiYsITGr0HNsdB3yrDqtQ+v3RVSR7ynTeGG25yVF2vUH1c0nnNIAkzzAGcMlaoeg8dZaDUV9
km5CgqorRgRdbIOh5miTdpa7TdKAMs1XvALoPZQ4jBtymGOI95VQQ2OANc8RCwLbUU5Jl5UOn9jX
JHJ1wBWAZn7kB/7C4fYTfgZmJLqXm8LzRsmh7WaxXHJEpDV869XwWZgGotnQJ4u79MSxtdm79133
gC+tdemnuhjGQvgqx9OnxusmUsGyCvLNUhM76di+Z6OWM/OTotfPtgaxUUiWkcRSTGfPuHzljJp9
6f8QwEvBPSqUB8hmyB0nYIALHsAAeG76XPWM/FIW1reIdxDHPPmfNjuLhEv72T47EonIx2S/LwGE
VQirB9LfT8SGXkTPSKQZCJ+DbKSg2Uc2nJg/aptIgJ6DlUERVIM20fxy7+UVYw5ZnYfghE5QVH6k
Vm0BZM1T4k3YSXIyaowl2H456w68+7GmS+0VfIAd0dBpG/B/gzAXxQpTBDLAgBWJnBXSFaQmdlO4
8r2FYx/sT5bL3S4VN/fVwFBGotK5ZoP6kVYr52tWOJOiSmfUM7fqLQjTEHo/ifazmCaOuhue5xTi
N0wRD7kRM4FHfGur/fh7OfFtx0rdZk/KQVnIElJzOiJX/HSH0kpZlK6BsUa+OQRY43RW/x/NHt1K
pY2tFl5/1hicoF4hd2lcRyH8PHopgTAbtm9n/l7gn8jv4AVC4mmeRUgsnI5PdqqUn4tWmZD/JwdY
TPXjIMmw/y8giPLgGgaLRsr2kwnhmbkMHuTk0WYQ72EJuj7tx4qXrR/9nYfPTDgw+JxavHqrv4zz
7ZC0Cg4+cmRU5/Mo1GJJhDkVFnF8WvdWU2pDkW1z886ETayXpzGSjpo6ms+DhwzO1yXR/ZJx8t0L
WBiGRwaI4LvnzSUPqv2qpmN48/YdZuxhE0gYkC6xk4aQDrW70PvvJSNbxyQDBvWgKP6Im86tlhxd
RiEft+r3/8bN39vJtapUc9WIwC5HRcSdXSFn1nUkeY9g8aZSKboLRL8OO6Oe4GYOBdWLzYEmKFX1
tm8r+T04FKWdh4mlEJftbjSNrAzoxR9+NuUUAXdGEomMkLBBX3A7JHz3txvpJSfdKudwCbcE6V/g
BQHNlNOA3FtV0lq2CGNQm6YQPacRg8nNlDYW3aWHJz/UHgkbeb7STosXzQ/PcT+333IICoiR61Ma
F4Fwp+IagnEqHT8hrSpKeBtqEDzFs/787fknQytPgoa2ZDgTF8Q0Mze0driqQJ/+XY9R+Cjvc5XU
568sDFxbYiqVx9WvQUGfzR9z4R87VuSfqG2jJABCn67gjC/S6vl1AzYfFL594v7Gq+KV0VHT3u2Q
ZdO7RJMGQUHM+9a22I8r/ihgQrKo9avwo6n5fiuWBFtwurjYtkzlsPKpENEXye2Qc21tehJ8AVPI
GrLj+wBnbQvHoxwhypKac9i6V1NgX6WgHsysxW+mtfCzlUJbt6ApnZgqXi3LzaIwj/+FcccY+H/R
xbDi9RQ5DJGEAP41+DAFOiCpWbY4A/KxFUGQtSlXHz3VB5m3ngCKwwW+0ZKex4M5x3y0NDFLZfRo
QENQzGBMFrEnnTBAsdh5Fw1MJ+u8d5tyR7P9Qw9Yun8SHGYot7KmXgHCw06IGw6YWg5oogqQLaZU
dXAq9sKA1O+kPu+rGed956Q9DPloe72nAS7QS5jVKuXpEK9QB2N4nV7m56OdBBktFcpc1YMvtzxD
1nJ9iKwcxlq44Jj82tUPbkNG8XV6i1Pn1b69nKcMLliCTaEUmxzUw5TJbQDp21ttK3uPnserfjyg
AhAFLpU0/kO9i4/zT/mfEYjPmx13cw/L1Xjc70b9VgcuvcnQYYkLhPdpp4WobTgkDKN6UotDPUm8
I8oCFUdb6mdJsSrMwUl5GyxgmjGZ1H1nFMCZnFpRhIfg/CSWwkMWsiWgJWTHTnpqvOEqgzQKztg7
0UqlJdQ8z4YvYsLCH5Wqd+8gXO+rrsExgHmk9ty+FoquoCyV0bw7iR6zUKcsEnfsoYpDwHj5SHOt
Qdn95ZYgaE2L7imAIBkdkesuebPEsXxgn3bGNMaQFLwNyw4y1kqjlr1vCjj/0JzHbC6WCLROsn2Q
/s5Gcac9RtY77uDpjJT0EucJSPdjie05jOy86kRyG8CzQUoEOfxGIbnEBWHUihqQbDtgTvtLEuhW
1QcMoscuwQk2UqFzt/19LIudBPK3ffB1WAxDv+gX9dMWiY/OQzM1dHFHb143Bvt9oOBdGadYwNbm
e9YccIopZRJSQ4xMW5lT7fEV7vDW+n9hRP9hkgNXbewBdVouhOnYJWXa6P6+QVfFMDnsJVhKbxrO
YgWqUz6/zqQqr80wKwHjTG/EXqbCS7SBo2zFXE6zOId9ZBeekNugXXRHulg+LORHHtRVr6avJxcH
pfD0akWUV5SmA5fPaPmZyBG9DsA6RNwIcRERbJHchD50tPqWBh19fOjNOvTzWAHjkSHhMvZIJ7rJ
YSozPf+OUx39wGXWGEFdodPx9R5JT8pEks9oR4/ZvYPaVv2uIC/B6mkYMdBeFgrXJSznF6bxZPU0
/vWd5S3xEdI525UFHEls+aVYY1WABkLDqTIxA/VkRzU7s/JXW+mBlDa/BD8MM2jvrxYJfUPaVmXN
0sMtgYpn9tcntVqNaEV++Vw44ivmHj7DELvVsp1guxsOpgS2rNXu7elvV5m//FBxt61Wh0NTsfIO
ecIZjkd8K35Bk1i1lBXXzQgaA0/hhUCNiMH5uKyw/C/31C5X3g6eKDpTI6rVgpyl3qkRCA1/MaAb
46M4XY0T+wKeOzlHUyD6CkHov7+lMwdDWGis7lK+6clNutrTlkTOQw3IBrw3IEt73dGXE52TFZav
LMoNEDzHEMvqJFsha874v5vBOlWS06WRaUu9m/cms3ryNSBYvzoMyEwPvdsWb/AcCPdmY9nqkRB3
cDshC8GdD+YD7XGdFNohterN0wAPJFtxGVj9mTByZ7ukddEctQBEpPQFqqVPBGLSTrOTJFK/7UaC
TPNK/4yv6jtjkzo4ODBuYkXhV6+gyY2ysNdz6v/qEIR+OAeHmLVEQ1WqdNb0GWWYjOmyhebP1v5H
+Z/yRWrx6tux9sEsMIDAfwgVw/tDKAE+7D2so0LeEMnFc3ezoaruiGVbJfBLft08Uz42B//3rMQe
E3TUb7ik1eRVOndsT7picz2C92OGqncSmUkImd1Be55OfMEGS995zPLHL0EtP3fi3sS1jeYYWXUP
Mc7GpVd8Sx7Z5bxs/4sadJ8R0a2RyxqxihqwY59+9KJQgBICEgJjXfImEnkHD3PThDXL9y5MA0MF
jbHwEEEmRXGpEABgbejN9hB7ZcNJaR2NzCqnCnx0RpR+LqHJntTwA4Ww0r+XKT2cyaEdRpjVBgQr
SBdvJhKDmEn10Y3F53CSbvCwHaaYZ+LhKnzMRaysLdCZK/7ieHoVONmEPP020iR4xVoeGLQSjlq/
2kEUDFIZ6T8gkT5+QGBdGYQIoBnFkDDMLHl38+0hPTtJtlzRvYWiFcf9I6jhtnqGcA86ARjiD5Q8
hY+FGdm9PrZ+fDhWVRjK3Nv8jJPPs2jupX/D9W2/aAYKBEzeEEWYC4En4mGyAVHgomt2g0k+hsa2
N+b76KL2p8E/QeWl4aWvUp7cDXO43EC3usJwuaLocjtcg6zKgAlwXxiTSDOatoa5f/FkdVOAEtHr
c6yGYSRNcnyfuIWrsWaiAjxvGiyY0+mFMG0++8UUNMVFqOVT+h9zcRNLQjU9pGNNqgLilrBdLmxm
1TJW1oJvP9lJUl6QK98lDlL0hIqs5TDbU6Ztp4+VgfW7eoFS0TINIuEKrKpAHhRf9L8XFm1Pt/kk
GhzSVFsSUPU3n8iW8GOYigR13gqPby5Mn+FGyD8ykGkJ9e7lkSik0qtwuo3nWLMzbr+0ioLid+j9
TKpr6FMrdVdiw6p7NHht81TSkrOv+vCpE6SAsytJslIsZXqUUW+2Dx+fYBybcfilaOJ/vnkge6xL
RU6NxO//HaYQFP0nJXWAt5k7ucbUZDcqtEtWQxX11Vadla2MvKrZGuItAyvByBEHk09hoxeDjFb8
oK0+S3LoAWMpYXc6oDPanh3QketB1Ml4WzqTSNj8elPx3gFY6AzMvZaY1Umn6ke1Q5sj/8tVB5RI
rPvmolnS38vVEHWdCYegopFZsilAacNBUTR7AAQVXKh0DrfNj6vgHtNfTOdhWov1I8ZUfYYlwAhL
piZVhxnNUdU0Esii84466VQbVXU5hLhP4Ha+V4L9UBhO5DJNipNS9Rc0lkI61FuzOGFd3NefrOse
Yq+0NWKKfwSJ5soBczOWM2sFeFKUT237VlIx2Vq9Cf9N6qdSNkIuVOO2scBbyKYYGu6zpQzRGpc/
jg8RM9v6Q1aDoyu3rX3WF7710PPB1TNtsHlKA1U9csZDjLfNE6pU18L6xwXTrHdpQyzPOwbdyaTD
9OfvaiKsh8Z5GjIFUJ08GTZoyQRzUd/cnBVegxxEss+E3aetFTcFQD2NU8n6x9F0dOLqkX8d7RH9
tpgy/2w4RmRchd/1PIvpluQT+fmfrvJt+xaQhAsnE5R4a8UgY7o6CQJsINJ+lEkPkoSbpJ/EgBCn
JknQDZxwZ9w9bUr6OyjDXa+e+y1GCysGRaPAXOA1YH5SJxKtT85lTPc0D+VJhK68LEJFSlDDIAbY
P47YkUJQp/62P9f4HSYxh427BFdw2CsHw4R1l+sTU79sSL2G0gJegCaQoZcLF6fZtztZ1h4Te7Zb
JeIiF8BD4iS4D6obVmpRUyrE4bBo7GZuFAP7ElWqKTXGhe1mqeO3WxRsc/iHcj8s1uZGMVM5KzgJ
xxtj6YWm7UEfPMunAzlmL/pn+cXfCmCb1ne5YF7UVgmSy/5eXXkIzejaAEYYeTAp7Rjws0+RxzkS
YNqgfwJjpOcadWmBYdtsSDZIxuE+HPe0z4uTTuM9DVDKZgzpGg9XRpiX/EjsXetzW7lSYPt6hCv/
GuqsrkwSOzUKcfi39QCn5RdcHedHELAwjySrZAySAFITWVX52EqydAkz0SrioW/cMfwX3lU/hMAe
Y+Oiw8US4KLDQy0A8OsBZENDKPJk8D0m7/B2avMEEHDlZGGK4aRKpw6KXCsTEHJO1u6BI6JSGbkX
OBprJorTU+Cdffkpodtt1/1067To8FCsaIzSmtr0a3UmS64x/X5bU0IVCUz3iePoK/dDb/eUlWUF
UXf/E5bA/1P6Oy0n7uRB8NDvmMjz0vPoL/Oe21WSiRwelBor5qTx2F9inTJ9pXlTC4v7A0NtqaAv
PTaaeGeP+4dnfGGrD/ISLjhhScOnhpUc8O89y75qfG0Mkn9lewLQzboNijuLyud1y5tBfsc20PQj
gA6T252iCiIzMpGW2uxb4mWHx6UdlRvP4T+9MzyZxmoVtFSEE1MByJLBvOQl7iNSwDcEm1UpuC6G
kUAywJe4TuF85motaLDRvaIf7/uOR0eJKk6IvmlSxuwJh3MdhsTuVK1JA9TAR6Z16zI61PqatOBv
XuccJIVUX+yuGgDvtwKPTusGvNozc/8JffSEMpKr1khQCiYlbu9Ag9IGdQW94E1dsFtu1tk0CxUd
ZNJFHCTAx5JerM86bev6/MQW7kNox/jAQ31MtA2L4g/gv9byPnWoP2fcjYffTKfgu+DzheFzQRaD
iG7ymbU+PpuJ34lE4927Y4UGUby5qVuDPbsjMi1gbv+IJ81EVBAfmqUdzd7bPL7MVcZ/+5c9bZ0H
0nxB5Y313xYXycU2S5T25WUuJR6yBSpz5krBD7NwbHw/sXcB+BQH7++yi66z2gVxFkHbFUfz2THT
5R+mpRAYM/A4EhV7+rIFRV+2t62ijBMxRmD1yhFY5Zh5WYJFBbOZt7wyVTbTAWBooS29g6khcZGe
C4xr2wIysNlUBRhpC3pZ7bq5iqTdP20hbOW4PP7U/+wkj+bQAfpPRBGch0UAWgoeiahGHkKZJcB2
0mS6dUgJgDvEG/NGbI57OsWz/h71hMP7xyYQGJET4KvRMfko7IxByx8daOvq9KIt2j+7tji/7SxC
xvFlI695EGijD5Cz68POJ7CO6xUlKVBHMNDqR3bLw7GaHVGxeZl/83dM2hZ4hP5uYvqB7S2cJ8SO
5xEwFy7/vNub6lC2y5z15AN7XTbeMI1n4O1VdQ4q0uqqgbc3Z9HorILWZfe0FeXvLdALwOlJngHX
Qvy0gMPGYsjzQRA3OyzQdXOxXcTvd4yRcQGsD/RL37qfNXwrHhnxygbVIYGrZbphLv7p9Er/JaZF
ceqr1MraoHC5gKzyGZg5YX/axbljNN2MfWRuJ4a9quAT6RGqJBkiVFMU7CmD5Vk3vZiCTJZgR0ki
ReNGE8i9nbsxEzfarLrpOhNJ862OJzmRat4d7qdz97PDSjmnxTKfkXnLJ6UW0kfsl4fyj9QqG2oe
tZU/ZWsfsKaVtxzHsI3gp/1cUjIvoW/jLmIjCAN/RmbclnEIR2rkZeEKYwq/RC8OFCooqzT0EkNH
8kAkqDdTs6UkhABLtrRgcgOqb31zv7CYoxUp6bbhY+2L+1aZNbUesZRssmzGMEwKxdf72T7BBsA4
fTiaFFIYTDpjWKqhqSlY/1nyK9MPA0QIMxgkFf3ij35Ydflu6ppp5iDxMGNiOD/v52iAjZItdsSw
vJkqu+7GO4mPxHVJlRAGXk4VR3M/08q4e4JWsnVSdXq1GTUtOxvKnwyE/nBBiOPWliseGCDYIvAn
HXbdcfB7/FrVqfSXLJDdBrR9PQWvHMi4VY+YG7ONi5nhenlJwug+qurKS+AbJKnBMKi77ttBdaGE
JiAuFcJHvmvavAGugw0DXgbm8EOKvImQpq39FzHkrhsCPkDR/xrXgj1aPbSUkcIyDBrCpMI7zSeE
x9mXX1Gng1gerTlr1pwLXBHM9PWDx1VX66Vwuc/hOQTV9FKpX4LZpQ9F9J6h0QjatIbTFpFFHTRE
J2kq6ggGVH8aU9ZeyRe85cwvym7fib/oiZqi955NV970JBAO54oj2EesazYChGs/dqN8ks/J2kVD
+8VFoB/T/64Ztx+eMjWPMw95jBqWpy2+6zRfCBNn833u+kDG2QtsMJ7ZgVS71WNcJ53MU8kTVwBK
ysXO2VQUuFp94YASrzZ63LwUtkuxSAho/vJmh7ifZaBXieM6vYhuDjMtfypg1teUwCJhGMtLvF9o
NyqdJjApE2qJ7nDtY2yhQ+rL24jhY7YuSdjXhH0imH2q3Rz00PWcqjENYGzxeGbTgoMNn39fRuhz
QYyVlpj1vWpGWzlb5h07KcYVaiKzG0X3S8EzfxkixcL2/Jgv27gM3m24U06YTRSuyKIo1oYA+tns
cbQimmQG+vxWfekfwTVudi+c24N/s2ADcNl2lmEVgLnNg7zr+xXfuhRX2K+z0vWv9E1p8BNU0Jkt
nrr5mad6MCB/QGU5A26/kGL7VNOU4vm6KhMGfpx9kiDjG2J7iriBfwYZmWpuaSZq2EChpqut6W+N
4sog8GsXb4sttvIOz0ciT2mZ2Pq4U2MaocLEz2zl5cs7W5sV3buNye0DDkVW85uGLJjL29tVanuG
sL92RTI6Pi8VTxAUaB7PkT50K3u27+Cuko171GYG5Wi+7y9FzknVd48yTV0IYMjPDQVThZ3obril
IusqBTm2A/FhPtvfSr+R8y61jmYJJ6DbbgoDTylPaCKitQqP3t5tUQmWhPKB7nK3611noJa1rM0O
1GtEiqCWmdHjO5FwRaNMJlShhYZpl6VnILbCqq3Ws7dixdCsCQ+vQJUirNYNx2KXhar+qVWtdfcN
hIS5bvhcJhVF7MkPucPGVM+UWBfkxjWQo3yAUHHDzKoAtAOEYgDfMtrtwZe5X3SRseB6bCyqj61y
2zRUGrxloEBN1R1toJTBhvMqwasUq3GZgfwNHa5OQ/kUC6rpRoZf51oHBuHiA4Z1NIjr9wFonOSQ
UYzvvOeH2Glu6VkCdkscxcFOU1DyWgxltz60EDFQbWhOjzQXX7lW8qmOxF2GkgyHGUxnLr4f0qAG
kHccdxRQ7J8euTpk6ZXOL9bsioJ1TXuHUBUXovpJwO9K3STvyKVWo2nuxOc29SzdGugPnJ2I72uJ
IfeUNHTqO0dKLn5yBWphwD2SFmL2YQhT8SgIfqOl3jAf/ZblLmgXXfNh+oMhGWsCT4Be/phA8jgA
c1s+j0D/D0F4KLbZdT0EfquUzogONcT3E2Ofqt4kN9N9XCFQzTrPg20THnlOnY3/XEznubTFBABd
Qq0JyUrMjYKDJ3ATjNL5i8ncjU5fIqN0dzEq7Xq+und5io/ecdvQMOcSHrpuMTwACM4U5AJSBK6V
+6i9gQDcfUNk8FAw5U+6Fr219j4a0FmmSGvzXz9geXtiBykmpWqb5jmPpw7I6PZoaoZBxeNhOIZr
PQOBQdtuFPtCR9ehujJxGM7C0DJLXmh45wykg9tks+JP+z+DXhd31jXEO33swVYd2dKXAw+i4cXJ
TzOcj/MHl4tzfg+Jv7RYf8I/7/XVfzMZedwHyqaYizHm4gJhI0iy/eERz3lEUfly8gpXMNg8/CRB
HahiOLrxiTWPjgFLUF3WAzWAhhbIkxYzPoWpktIONFHUyTABR8+Pgnyd0QnFUP64cmxWxlGMlWya
GB2tolVu7c4y7b2FFYarpviTayGsYAwKt++SuyLHLAOAhl3eUtUzvtW0IOajvN+Enal/dWyi6YU+
Nf1Z3Tdfi3yDHxCQuzoFYbGVEFg5t+L+IQ1AUJi9fM86RFArY+/Ra/GdW1pkHnvRIkmzQ54DgNwq
yF2/cddIT9McuM/QY7iqMpQ7uW4e2voGsil1bGihBaaOvbmIXm0TNdkAxRJUtCtCxpUVveGXJpao
PJ40ClcQt1Pu6WhGtqm55G7R/9RY3mfRP2pEAAkdO8ABxh/YFFyzxgi+MOdFjo6pwGJXcFiWWOVT
XU4KhdAonOL38LLsvEW4zAfkJwcGsQE/HgeUu0HG7Mxdu2xIvpCylklC/BbuXZcWdrDnP+AWBJYP
pGViQLh+dAyLVYyvtH6Rn9rk5TXQNJjhQnG9X/5Vvtta86BUv76z/Vi46KUopRyWAm8IXtWa7Ziz
5NMEt6a5UvfAAgDPTKMePz85Kqg4deDClOglmj+lJz90WnmETSCfjeA/rsoRlaAnb9t8z/T3oan6
Hrvm/n1YbnaHKePyKzT0C1nAvUDB1Q754IzSWLS52P8ul7TdmTyfq5E5dSkM3xgpy8syvRIJDyTT
0e0qtqaBoZlw7wkacB2zaEGomqBo5Vd1gR1nIGSFPpQTbdDOVBhaJxPz3Pk6D7EyCHWNDu+Bqaqd
ea8sWQ+uzdBBNrI1v9KExAdDB3PL72jrJT+WTnB5aZP945k/UWrJOaFiFYPK2XTdiYbUSrk4HnDA
ZuPjE5A7P6iluOe9mn4MTOZiVUX0BQbwgjHFflPNmgR092gZFqWdr13K5BCHN0WlzI1ocVSAEV5K
q47i/4UsJlWEM2ZiOnhvPpwVqRNGJGgeyfeMkOOgzku5zeDBmrY6ylehxdDlk9caYzSx5z5O9i9T
x3FIRQEiB+cReYf+A+ZCxz2YpLcUoF3zXjSHxPzAPNNyklFA4eJ54sCml6NWpdxiXX+6TKmMMpvv
w3yRP7aU8MVNJzijAAN2gn1yE18h0L+o9WSugzLq0q+xRtaMg2fUC6tPdXFB/wjntD82W6GVd1Pa
/hOxuWcFiuXi43KHSfIjY2mADXrYyGYv2vozdnrpfAzNGrFUxeN+0dQ3hy02QeFLHbOCV0Ij9ZQT
/h42QrIOjkDuhzMvP8IUqa3gTZmjIC5IdDze+oeR05PF4jmkLq8lawC5e7xXPbyNiJJ4P1ENKnRF
8AQIOMcWb96ghPfB7SmwwqaBNIXEb/S/SZSW516GPSyacz/cbCNhthE3HTzsUAhox3x1tlq7uLFf
GP2YjuEe1Ez3Gs38uhuIMtmo4IfJcWXDVHYCemiYqJgoAx7R/u31E4CwRdWGkO85IXyUSP9RRm3B
5m5VzZRDZZa7V/ZK/QnSYZWg6HbPhdKvdm6ZW2mCRffNZcumkprzKDaRBLKtUaVuoDa8N15TZ1Qi
Wk8YNcY4aeaVzEJ3xpLwwBmdJ77FhOqnmQqlX/8QhlAz/lgaL5Z3d/qBd7+0o2A0zwZwgMLw5pI8
FAz3JCFyTx0uDq0mxZHoX4cEidTpdNKLXdcQEUGpVVW8vcH3ltpw45fvRpyCnWCBX72knH1G610M
MOjLiGPv94OCNnHZS6bskjWs7WPZRa8RhrVT0yXutIe5TFAJdjvCgxk4i/Nh4GzR+wGXdg2uEXZb
cfH5JFvU+mfjpx+JVo+qWI710qRPNVV0Ty/GGHXYPfxBWMw6dv1G2Q7cWkmZzeVQHoAmcPaouxYg
X8ABNlnaoiuggT1EiQK8fJMxBsP9GYExmacv5eiSqNRrFSHWNFyq0pPfcB/hFjH7ADpZ1+vDVYpe
40zTzwk853QtxWgjGYieLjKyucNhP32n0eVo9h9EiMmRAFv5om6kfa71aToO3j9/r3hSlyBGrEUS
bL41nVtJf6wl61TdhnEM223Gj8aGks+xTitvEmAB+PtK2oWMmNET69ShiGp0J53AzjwWWT9nM+70
7HcSBP3GuUoqlb+ycnUQvwu9NTpiU/DRpl30i/d98/fv1aXGcx3+MgPamHVzDRVUwG5j9mXvlfwx
jsA/bYEYCCs2DE18DyW/VIHN795sJ5CLbbB5yKudWZk5lU2xcBPKCck+2PkIC+zOR6NFb9z8HgYd
k+tE6tYPFzEnUgoJTcR+rTsJdG+SiWK5/zkmRCMnx06fhIuf8uIuWWH4TQ0sKZm4lnuoz2BIfpW4
zaoQeKt/NeIIDl5MoyrAVxqjKAKYl51WT7L7SDeKpUZsnNj+j4lbWZgumsJzr/YBIj1Bc0GUKMq/
FfVAx4f3DFdwUAs5R4h9CRa9q9XcC6XW1ZIlbo7c1xTmZ5l4vnteIAuLMSkTz2E/Svvj/1gRA5WF
p0QTWG4oDlk8FydJn6vUlhCXDLdNWOS6nNToXa4sbO1OxsUX1zK34B7KDv2MO1708c5f7ewM9ziC
mmVQT+WgHIVvJV8JOUgGuhR/K8/rNkDaD57YN7UOfYbfsggU2NqH2A4Wq5sGezBojpM49/8JsxIq
6M4d743rNYzB6m1wzGaL3Ky5EWUrigEYpeWonbdExMD+0uZRgPw9zB9/SmqUErISB8QV4S5quvtY
reUxpvvLyySwxxKm1p7H9Hpi7A6GDa+5QY2F0b7geQnHwHz1vG15rtbwrp7nl1Julr/EZw79e8Cb
dS46LTHMpc+LoNgkur2FhJBj8Y/wB+kS1m/Mu4tg+6Zb/gvPQ/+h9RywwjTYr7hXfKCwSn37GtPl
hw9zexL5cQCxDz3xfNfTUdsSzx5CK2vRfuIsAJr+Q+3mWr4mjtS3pB/UwbXrxRCvcjUvk0H+Tqjo
uXnFSvs+mprsc+Y/0UVpxXM7OofjMv5GWgGP+xZWKeuJxw/MV0e9LQTawSrWLscX2KR7WTFQztTB
JuxVclHJsvQGx9FDJeaXWhve02rgYxwxTSPsCYpr9Y/yBsrl6sq9Xe0DSmyhRKC3O3Rg6VI8qN+m
5iVY6HfDmelfLlE2eZ9ZL9zw8YtsxPbi7K0DdNCDmmr4L3x+w5XIp6jiprD5aan1H0593w6jrIAU
HOBKCREGo1XhJue1BptGt1x+lj/l6zsGlUJ4AQ0tRw85LVbVHWGwNjpzrPPYMoNmqkqvtPCTWhWf
F4E62D5P6+nVfV0f6SBnWT8I0SuvgGiqARAAUZzJhjpyxCfeortfLq5pWtjQA0pDEv4+zZLPKpoA
I8rZYqGduPz4qfCZL0fbOMCOu6cGja1v8oWMpVk11vJYRd1WQgxEpAjs7B9Td7YGrzEdDjAlF4gc
p0IFDY2YZUG/Tc+AYzzFMVSFls4OLCthzzrx0tBQ+x2GctHGeeapSJbBlAcw5kRlsjCfIXAXeL51
/4DNqDgpEkKv4CrPC24oKy8XxBTZqA/8dNB5alw98Bgd5TeIH7oxA7B0U2KAD+JqYSed9Nsdx1Cg
3MaYJ4FZ3qsZMGqN9fwwwRu9ClKk0HLLVcVH3ulGOUwXSEm63cvZdUSEK/KCGC+zxowsqKbq0u7+
aANqOj+HOuIcyGva4vIFBD1wT4kcO13LBnaNuJzaVur1J5DCRmqmf3WHvyom9PuVscLHO4rLV2+t
IDTVlJjZGf2luUrJtr7CUQY3xMGtO7MM0+3wQgHTLDs3d1r4mGD5XBQgkjD+MjBS8+in8XrtP+Hp
07aC0FcInf9Hg2egEnEujdmNQewo+CbYWyYH8/3Yia32p3tp7SwpZP/fj2IyZuK/lel27MG2oBXq
AczXjyaClVdVqhEY6m+DA+8WyM+LhmXmsij3u519AZwOPo3cbGHL3Nn/rqCS35IVDxqwJJ4o5NOo
Wzrd6hCVIDTLZ4Xl/eGRtBsrNVgW0rjTKlFeYdpcXNd2w+7afAVjpdfVObL9S+zJhzMgRJ7QXUll
nGT39mPQqVgdRlt/Rc9N1g/iZJbpXCQbPLhkJzFjtTYoDfBRGI3gVbPH6XBzbgMGKhPPOxW++Npw
OsDSePT24g/vtgvXkMwC1+2xiyGA0cfvuUBj+hCkll8rJBXgGQK8la8/HP9fBidPme4ry6NrSCcr
O+NAsj5z5GAYzn33npKTW1buYbeMEaGF28c8eEk6Mpruqry6FaVtUIcJmEA3UvwqXGWWTYFI1rFn
fSfrsIAdibd6easgrv3tiMCNwVdi5mBJSTeHYjV3rOrP1c6uUeDrPW2YEe7xjnGf5GjDU8mlUPq+
oBWziguzW84FS58A7zpyAe0TINF9WSDERa4eJ69IoNXFRTLZ1GouoUzKg4z36O5zk+kSu8xIy7VV
lv5KI1hmXwkFyxM6ueMS6R01/RVudtnmyWxjfBZZWpjs9wa9qiI5gQ3lhZ3mUbPX+md9mhXbWcQs
qn1QAQ46u3GfjPDEK+GKGAKz6QW6HJgT9QKsk1Bxw9/l4D5/cSHC9i9TICENdVbyqUjIrTctvxjE
Tm9Q2bsH4klhvybBUE8sxtKKWDyi2RuvDGiYcC2KJrf9B14AdXxRrrNim85YZdJRbuCl1yok9Ye0
OaxwFUwMBKFwfPrGM48ZwhPQNFRhk7QgNDqMfC8wh3GDeETneohRYRqZ8CpBjwQPHMJXQ4FmwhsB
8pHW7QF0uIZwm1/3ASVIGR+SHx0FA4zmvHQ0PtQqDNUENZw5rWJzzITVckXZGNZ9jZPJLqSWSo3I
3noF89j3FEuEMXY0ARhlP9bVaGBoMxX/T64Lf7febV+hjuW61ssQ14MxoPVyC0yeJRxLUIQbG/Yv
0gzdDvMRfFd/L9lVgzLB1SKTndb4LfKbgNP8pMWzVBSiOTZL3vNHiZMTOPa2hINShGFkMJqtW22P
d8yyolJsQK8ZeXVf5e8BkmqYeuQsy2tdhK6x1P04fclboGBGAhdcnWIUQUwPDujly6J6bZV+ZQOh
KYDAQPEgwuZVraM9AbYAd4Deu2vo1wxkeSrKigb+ex/S13cP1hiB2IOOvqee0imoOtlOfco1qBfa
3DT1znrhiFEyklhu4972A39Lywi7aaoQQgYMxQTFG+pmXqH+uIV5ezSSqt6lpCfMZgh92BjKyDnA
+SxWtpceyXWbX2Djl2BDlZ5gLJo2UDRVlHdtIBWyu91UJmDjCgX4ZOuLeuMkELJvkUE2i4Y+aOvh
rGlxww6Xjf/KmY/asT1Tscd6xeOF5UKOowRdNCW412ZKdbRfXqMzbP8fOtetnPs+txIb1Me9O1OA
huKpVnjU57xoCh22EzsmNe0Kj/nEr1yIMFyHAfMSDv0afPZgXoZkG5SAhVb080G/hOpi6oVTjVQA
ugGzJDtSL//DaB/PSfxzH7wDtSxY0arH/+x7CJT1guMoYD/C792b3aLD1kmXQg8vQ22j1tUM5qmA
mXr7jTARSOzPJUKdAwTwOyoj4qLc0An+B0H8vJmhk19CJCvs9/2CEUmcXeO9NUV8LmVWixV+eLub
DfM5OsFFMLHmxEr1ngQp1mGicNaBjN4uERQjeVqfsuQnquI1kItaH9/TsdisxNJx6MU8XuL5hgeq
TPhg1zCVUJuYgzQa020FCM9Ex4sOYayHuQzUC45eIWISVFOJ2Mbl9rTfQqdx20oNt74FABxVM1qH
fxn7J/rMYngJAGiddDxaOG3a5zT6iyJdU3iC1d+bHK0h1QFbVV19Fxnze4ks0LVTkYghdQOL3bYD
k46vVpvtsBlJYYf1bhNOMGz2bcn/I65wjHYX0HkHajjy2J2Uw2gmDEwZqa/tPEUC2i83XHb72X+b
mbuR4wAujebq8euqP2o/5WidtSfPYFShOYjbGhHNjw6UKBn/SndxiB+MSYn/QQkotThB193a/M9t
ANTcn8jcwczQpcZ5PDGiS2lheE/wCmWqbbe9fqXBIbWWfKMDrb4oFGlIb8SvfPZbfw8Gq9oKqXoh
vNWPHVLl7Ug53PPHRVxHZkZhFhGydxI9e5nnrBUT1/msHNp/6Ixt+ZOybNYW3khuqNrl/oLP/gRF
HQKX2U1l6LHmRGF3zESq1bFdslMqg8zw82O3f3be5Ejl6cV0PX1VZAuXVz2Q8GuB5u2FvcX8DyFv
oRto2q2YUGs6x+MUORxa71KVSBEHg6tRvKi7OBRujVtml8RHVqRzgdxDa8ORJ93BA9McY8PSrN5W
uQEAUG3PreWmMAZimoZXvmW6KfxB9RZs1Kpeze4m4J+8uQVsJPBM0Xbdm/Xy5FpmNkr43DDkGNAF
FyIRbdH11hASuN7rZPEzkn4lQr1vlegyhL6O6AV8/c4Tv7GPaff3wWSulTEM/WRC1Hp6+FZwmUbM
IWXjClXLN4vtejMrLGVNkYUSY5mYWjGY3acxSwx6Y3S3P/a5DZwINN2jYVLTCOGshdObLhsqPVMP
pnHYWC0anrwoNObj1pj3JhsWoRtBPGF7g1t6yvQkD5z6gUHWo1ntTnn57EacPwtd0jt9PiwKPeb6
QUNTS6UXFvc73n6J6qP4xdPmIJP9iHQ5qA3WeTbrn0Hcirmc/f9lqnelWa70NdGWho4mYZGwgo+4
u1i/Nq3+dRMlvoxm7fs5ij3wXiJfrN+QPRtO37eLobFvT2/koELvBZvak4EXZnJoCsacNjT3bd/m
iJiN/1QpmkeNynQuiBzSbqKC33EomcV+Fz9INjNFkDeCoezDUHkhs289uDru7bqm3pDJAICOewAE
5l4kAqQ50tsI6kr0n6saE8gfcdsxTzUc901Hc+0bJxT/h9mxFiqEC8xjuXIxzwGvp7CuXFt2EnWH
ezHaDEeNzttn3vRyESOvMNoLH6tDALsrUoPdhjP4wsV59rA413S+KWhSjZWDzUx2GuSrw5v8043O
2ohXgemKS2TWZohmjSNpNXelSUv7swQ13CNhHk+ZLtlTZogh8yZLRWcqogH0lKRCck0Ok+3S9CW6
d3Rpy9W4MgD+URPC++PhzvXd3FVnnRYcPBWmCdQJq4hL+XVhyfCwvhpSDUgxqksuTh6JEr9iq3E6
D8c+TcZUalMzrtTEEi3kq7qTltAz8JUnCG1eRnXC8POrLCYRXZ5EzflK+UL+eif93nQzB1O9gUgH
T2YBFvL29FvY9mneZPhgaKAWLTVWECkW2vJLJQRAzO9UGNVuuJcYXTbk/EWKuqUdlV9uMVV07uAz
+c+rQMksffWQNtoLmXjTXC3+lLakPoAFJcRQ2i1NyZGlCQOd3jtGvdeCi+WA7/eGC8fvyIwj24Ak
l5YVA8DHUEriNyKbFssXr255P2rYCy/KQJNLwOK0oP52CTbA3dyjrbQTNJbW9F+H/YAHbV560u7V
zXcChzLJMjH28Tclv9f17IGZtYoPHJAn1szzqPyWJ5HmHj4u++Fp9wrLw98BGiDzgH06EZ9kQyq7
gOW4RPYyfFPJc1T03SSys9zADa2cr4fLncdU9KfsxASJmfskDzM2r0reO4C9rHuhsDpi/31bE8Ca
l6bMquOUgE8r+GEcMBLUmZWbPZFQ7oqQjkBhPhUlV2uPYwbygpv53y0NXQCbbSbRBNQUjp7xwvzm
Fgke0Nc4SnOupnzoxAAV+PbU4VkAoLLHYefKXUaIp1sjsXMbn/iOgU4nivSGkOqmxcO3ivFRJ9PG
GHQ5JWnPQsmU0Y8mxjKOxHwng3e8BEygdE1W4jVLbgmG7InQqk21jrdeRDx1QMrdZu3ci0MWzacG
c4wARO9WNUyGn62HKJ77cbym5MtHW1lZGN4SQiKiAPlsFJuVw1qtLAxNXhU72IR8t4A1kN+yuYlC
1b3aFCSrXzZHwkYk8jIdmURK+8Xv1P4oU5Q0c6tCZX4OC52WzFv06gnHoTLJOOFddtUKuxtSW1FL
K+xln3ZyQ60rurfituIJpsakOmPIuxKjmvm+RMGf4AMb5NHyiU6cghavFaZVvYtRwUnwtW3QfoJf
Voise7AQ3kl1pXCTOIK+8zFHDQ76YdUxBU4H2u5Yjdd9EbHwdGJ5raAmqrFApNiPUcG7Q2ksTJ8j
u9iW2L1108tgkfUuEsvTOo7C+X115ieauw/Jl0AXZwS2FiJhnIMUe+IOTwl/kKuVHS6E2i9+RRFl
dDAmJIMS1AOphqPt/l8Nc4Kq9IsQMv1IVFH62VyPKv9OSiXTqoH9UYjqyoXd9bHtreWxK3YXVtZE
whg9qTYIoEIsFeWCEsApWxPNJ7j4dAr6V9iQuCcd6hi+3M21OsgA9Q4cKd1mfnzWbHXrpaYKf78n
c04vlgkoG7BrnN8rMATNMq1VkyiPNBH3wmYJ76wKeIf5VjcPZXmfhVAeKZJTYd8TF5JvRcafIROX
EXCOLmS/1adokglvIHXPHae142OE64C778tKOV4twOOMZcvo2wOcTpbAgMo/pOHHGPJ87PUeNEXA
Dlx+fJ85SkEV0PEDQAl1dzrQ418DjJoShoeqfa6ZV+iN6RaGifxXkdJACwn34rp/v0RT7dpCRqa5
YsAh4Zma4zX1bmpxJ8ikR2zkRyN3PBwPBigkuIgVjMufTdG6BeHCV86TGlGE+oqJFqkTxNHsQbTh
FFsmWpLPm/7WTYkxb1UdDTZq9/Oo6KhuHJBJD6iIbGdO1DNgkcq1sQ+A66us/qw6lZw8dMMmPDC/
32XMQ//SJIK9Edu5eTph19gyWP8mr2HR/1vnRxCV6Asnkx18i70G/5hUiHJL5rSlo31HHjUg4Mrl
4oUTHLGqEpADZF3CzAHVCy33YtYlnawY1+UOU/Z0q7aQ1aU45c9VPefTnjK02kjC7WeXTI2O7Jk3
ZhDGnZnkLI7JKZOmR8/VH9u6gNPQAqzy+40BIYQmDyOOZ+qR9XzhTHnO9+fZWzeUHRkRHZtlJ0pG
Tq8oZYWhPgo96V6vj/tlcmxHAlVy6V/tNSHaQLuYdKD1IMxMEYi9YLuDt5QyXi63bmwgc+q6Qkq8
hQxO397eA+1toPcVPGNgVTvTnceLdmTq3Zm7HHQ4Fob1M3ZrMlaTgM/UK/SAPV6HkHr2x0Z6qxtB
bmy9hFwZLQKTHL2V9ar28+B3zVi5OpsT+X1Ya/CiEfgaYtcpWiJp8za2VqMCaQ73VPzpmk5IlwFJ
HFeMfrAubvIw/3ijzQLn4S+OkA09I/kBtImfc9axgDahqiPuXEZ3KkXGYwJL24onLR9o3Iwtopo+
oeMBdgSaMsgbQ+jSNO07OJS/A9aAYctxzkOhTvlN01IJ8P8ZyBbbTzD5usSU49VR6IC5qc9t0Be4
53fXFMkhPo9BNIoLp8Yb+hi2qZBDsQQueSEfx/X+G8+tmCHBRInm9Pr8fEG4pyzZx4sJhYh1g/HK
bMWSomYeNySdo22J+WgAO2wy0by4t71xBGfMGsAVPNMixMCg5+QmXK2xlvdq3ZRGrngQC2CYm6XE
kwhIrKdCQYSHxMfd/qG6DFQsM/fYVRcb+nUW8MjG4c0mWmqvHxVuGUMCrhNkUR8CjHJTYbLhW5gI
RzTlA35SL++HnRGEXp3YIAIUWHhaHXI2ioH7sKxfsdTQuisRxWJY+WI925Kdnp5rE6ehHNNCh7ZA
LT22VBD10hlKfFXx4fljAuQkK1q5MEHV4bhmyFUItImllzTqvN79T2V25OKAUFV7TyL/C4WI7WCD
ZN0TVBbLAJUnrNpG92nr3JKF0ozwYNXga8yt5vBA4ZjMx+5f6PZ/TZnho3+qHa9XKn8CmpR0EP7y
bjEhqtDKihOa3NnCXn62auWa8GSK5CgxtuIZkzSVmPpjS0rYnLxICUDNH6CV+bIAjeGv4CTFXHb+
rRgH+JnG9V4qu28LU8A9YN558l5NWkos3yXXv4fydF01B4QVqpCmBQzQxCvcASHlEY9QM1MnU98A
B5KR0VFR7kzHoVBwEOG6FVfN9tB7xbKCbLbqvcdfLk5fu+4mLykvG0jYnnpGLeeMknTqGwYSDC41
TYulS8WvApslfW4zQFtEB7n4gIPxOvYR7C+0lU8045Zug309A5Fofd7XwK8lDR2bStRXRiX7BVp5
iZCrAoj5EDY2lX9KJK7qvPZGIQGMfn8diPeDCnCDgOB6XVqvnwgFGB8N7vIJ6eBEOJy/OMtU7CaR
hWkcqF7de9tPLfHKM/XlixKldu18BA3PKqHqoxjz5oh6pv8Gam3ANx96kvn7mOmzjGpPd+80S+vd
jWA1rI9X5eXcWxO5OexJyEJ2oTvxaVHd2B48qiuIbMHn/s4MDK3xHCMLuagYb1mZChHYoz133wbl
kzAlfE019fWzQnYy1aLSjZz7CqLZFYVXpG8+2OEz6DnTypRYlZUtoJ3pN3W2UMYlsoyh3kVPA9Xq
kW/2B1FiZfnfcUDpAa8kGLiuWQ+658ab1BNBAVSsakoU5VQnK0JN3QQY0fmzN6ndnQEeGCsejhxn
a98fy9KRJ6VrwRAg7jraxOWK0d3ZgDpa+isseXY0Q+hiVlzvI5zewdnuclNq36GdH7fb5oQdwbjo
hUaW+IMeI0jpBcwmgc0qJ/qQAkHIhQMKKSzQI1JoF8gO9t46NhNgcKazxGRU4VpqZIW2q3S/OUTO
O8JvE6IRs1tCf/k/XOGLuuGHRExzq+4FtRNNN7O6LHMzyumbPLRENeLI8N9Z62dhjdb3ZFPowdRn
94sRbc+WyfEmlgqfUzAhEANOiSptpJ/wq2gfk/Ttl9PAyVFtRdfnzVcjmx7vFBOqwkIxU4yQG422
kLC+/GAAYdsHqDxuoO0Y8604lCL5iSVXZ52GWTegIAjNg2ByW+haCSU5e3AMoJyKrNTpqfMB+Kaw
Dvb7t6glIitpQcpaI8Jl43bKv+oiDCKsThDBbISdzAtx2sac5X/8lsu6Ns3dgNJgJdHyPHe4KjOX
aqqymC5nUuonKD6Z2n8K6Mz+F7XMAr1z9NsnmQB4K1OcI8L7LiezYcTnTugbwm495UmsfYqPQn2f
R/5hT/mlu/mn8pjKZN+vPKUtH+fFEY4Fmy+ClMGvNNCXWIOzYEvVv9tzfrR1QDMhRXfNPQPhg0qK
SJwBDBT7/qlILGBFP4yvnSBq78XuDGp/WzWtLMeZaa/lA3VVYRp2wy0C5w67T8qunRsTeZajIhc2
bOfbhFMApEq2nB/YJBnk+zHivdBLo73jW45H6RuCxN3KkR8Hy6Jg72Yc4Sq4iQLt/5ElFNJIhFVe
lv+1zRSKKcjQuMII7nYv7RrOs2/M3MUdCaQYJE4wuRQD/wkbHYG3y4Roasrb1TGz9BGgnSzzCLrH
maKljlDlrn97MwMjsJiwUB8zJYLYku0jGOPDG+yimYNmFRq78pCgHqczXz8giuCCypYmVdPnY1k0
YFrZJDYIaf9XYKNO1U1Ya0rxjuMcLoKe4EDrvsZx1MniQLG+doMHcw4Re2QPm6cu6jTLkdTTanID
sE5/rRnwuiquXgJ7WJIZB5mbyPUxBCY83hCpCk86aLHoGJD/DI4dsnNHcb6ZNQsnR0wsewLwKh2c
uRNPtmadz3FTqhJxIk9BFYqjO56ZLKuOxCyJ7Fz6ZbIZ3QWzjkUAZwqL9nTG1vrz5uqQazVZThLr
SsgcnzPQLLts3yk1qctrwPWVb6CExIhzTkdAh/ZWLkXmNx1I6LHqU+jWJ5SnaYq0489uc3ObDKU7
6HWgBGR51ER7YLSqAGhtocwbSBf3WNfM+A/Bq/5SRGWiCK7EzKJiJ762gbevgfGM48KlfOXA4dEM
wOFUO9LzTZcocUgN7tay8T4NlZ+ZLiMTiyXyCnG6ckd1UDLXZZhOoyU9i++h+jFbEReAgfLiYghW
LdV1B8jUdRshI2Mn1U9YklyOgJrbOc7ghY+KbVaEBREAwVA5cXSgMHaeer2wQzZ7s4f5LfFBFOXL
8EWtZgRtV2Z1sQtn40hrrDsxh9znhPIPk46YPTM70qnmXuXuXSJFAq4jDsyobvQKAx6SkHGq03+2
ythd21sbxT72sq4OQAMMrx+ly6j+iM21pXk85vX4aAyN8TjrZ1NRieJbKtNEehi3U3K/NCnqeXyR
GVyPiCkc4QtPXXzrDtMvxjq6boo2ZmfQjxo86dBLFWa2NYa5HxY5JXTA9PDsEC+cTlMyseQgP6Uc
2O6qd5wm1XKK9NL8N5sIsVKdT/P2WNmpCRGjaoomdUixvM7RPRwHWNTF+RunXv3UPj9ZywR0Odok
1YQTbAja3OBNCIHTVsYAWRUjDQcLD0NhlAAsA9whBYSQaVCA5bf8Be2hQh/j4f8g6M9dx1v0x70e
FS2dmkqerTgRujN2e9hDaAdvIJmJDs+HVx/OcFOQ+NZg5U7Q/Q1j1Ew7cUbiTKR6Lqxul4Kw0CbM
l5aC0tFgbWK5FEbsVZrZAJPH+B7ukz4y6rlo7rDD8x5LogHYFrew4j1zDqnXr93yrC5Ii111+76S
JgYVtvIQzRTMzwL7LagAgqPGlxxVlWyeGlp+6QQc22gM6zVOTHgVuLa/6AsjKj+xnci/vd+SBJSJ
9EQC0LLOtfppb6JfDRf/fFNbgM9Agn3uo/pKqwrOAthM9c0dlvP5wpd1ufbzD6hGlEA0n/58rGLj
iCq7W1Vm7RAWxOZNc5ZvOmRAMUe2U+ngZRnookIdr1Yqp1PMeHDmWTwchDMg+daYl7XRoV0wcPkq
QQi6BSqnVxo3PrJBx9A2ffy3Pn1vWSyiic7iP2PyCVrA0YMpATqjTfWPElDaLUxozr4dDJ5gsGE7
DMVt0m0Aeicec90XYLYg+fece1SYSkQwC81oDNGRWEjnivz1BrGzczR4M8Feratuv9QBEaRXOAbO
3DQTJpuTz5A/xA9CWiYzQ80uW0bncaURe795G0wItduYbujUwyb1u7abmeFtyVGoPWPMDBnYeUre
7O0xWfeQp1xRe0LpqaX7Morw9XZAVPSAsXU4XikSxNg57TuEcb5x075/Dky5rmOOW+t5tBCW5bwr
A/GOE67SmHo+6Mu47lZty3Lqj79sOUChLUIuKKT4kSamk1KNFbOkRVQzykzwdH/7PYO3mLJeewSS
kUXAwOc9VMY94LwcadcXomllcci82TQgQ9zn93GSBXu4LtWLzsovFnBCWdeGYEAdtfTFaLflpCK9
a53Pd7X0u2rFc5M4Z+VyA1rbEdG801cTT+tKElIwZ5FJ2wL3VwdgZXcMgb1DxlKK+7NVlMcYw1J2
/VRawz31MbEBJba2tZTQC6qh4QVjBMhcV9BR2vM+InXK6zFXEjl+9ewLBpI4CA9L5qmPyNoyff/4
5roziISZMOR7xAJ7toJ5mlHG1cVemiw/V/5n8vRRigSaipSMm9ThgMOZbzTBYgX4WVnzXWFWcUU7
pKPexNJebRzP9h7fPxUzEQ5ee86VtpYc0NZd9tSK3DCOZWSE5t0VF25AgnPkpNOZIG2iNtBWs4aX
tdl7zb6H9JLkx9glFccXUiDoD9qxduD7WJLtOWMTWHGT3z1Mxr6ALGJG3VgzXpwcyBzNFGIpoYTF
/q8E7o066E97U8y91mykVlBQSXNnfh949/PbiUNQ4AjBry4yj1qDsjTXc657GIQNx/gS3UWayGxQ
+XKZp3PYkMXSCypy9uwDReXtbIQwEe9GbIcaQc+tQIzetF6hK9KDmSRNeKNiXraUaozWXl0R+IYH
XkvBGk68ZDxjLNLOJSLPTomqCY0DQDoQg4e587sC22fNiKyAn/DHfpI+ee3dX/Aj7dRDxGKxzKBH
+FNiggb93uYs0ZjMX9qZbVOnGI5HbtifhUP9GoKuRx8YVSVEquDrLRJpmwR2y3BOSBJ5JM04zpuz
NAXqhfDcy5SWWr2e8yX0K1kot6KwjSpwg9PMwQAq3tyM/ZhhjXA2dIjAkUHeByRyOgjz8hamJSjv
9XoeNMtYMTQo0s0yZGIkBQcwS1wtnTO1qkuxB23cMdt7PpFtXqp7fRg7mXHPmllFLVx7p1N0gbG8
7yn28754iUoDWbnhreTqEVXnPNtIhsPOLVULFB7/TsZgNawIyMz8JBCbtT4joJhbQ7YMaxEODtsI
9F5yuqcNWkcEUjwN1stROqofzQcuRdjXPs9uqjtzuBWz4JlYFimW+a1J90n34X0hkjoPuuKHQ+AW
XpYg2bL987YdB7GSdERJw0g3cVHbUH62FE2tHKL4xlcyzx/5TfFjOo4Zxk5kaPa3O+nmSuoNDssk
ULvvUuThf27m2ugxohWC3LwXU1GKhyFqxrztqsM9rXN3qP3eAouhySf5gsxMbEfJXevN1QV8Vc/i
v9BbsuVycBcK9hgO1PL8g4W7hlnveLw3igimNL2MKgemCiTlGWBhn9/dNz6WhoMt6df3ZRyzUvvG
e8EAxFwthgBn9/X7OW/IHkii1jrry6BUL5+jqGCEopr3VkVrmesfDyrhw1f3zWU3PanG1BvrYCQ+
e7Bx0wuLD9R0X/Vol9Ou3jEe/vpUP6V3DCo8rPN641wZ3aX8oMZCvjLa/PQQnn347ealOPSqj+Bw
nqBGMRzbWkX72FTy4FUXvgHObPXRKC7rhA0gmKlLG0JLavVcTkm+B0ovdRy9G/yfBKsp5YW0I/tx
HzRgjkWgphtjDhl6qLREFSJuYweVetXi1j8K7WOmaizOLdUx4L1GXS1CDzVHvvlQb+mXYqXYxu5Y
pphTxKF8Ckr13K8oq5+8kdsl/TRj591oL2QyPUx+6wxoV2Q8szgqiO8gd1NEZ6pU0hdkhRC6Zreh
xvVc01k11IUH7ahM25johGpbHRgOzhrqXrp1dfQ31NVMA4NP6WANZ9DYBIHtxdOF3SgRUORKndEz
qnB8ie12dvCwg55xjGcsKva1j/nS1FxwUZWbJLE0D8/UgrcnyHHP5D2gLvGTnfWGxACNYxJLgYmP
aOp+AyJwaZEEukiaL4m1KHCD6ns3Zoopiv0pjj0Hw2vqh+8/LptIQ1kaFVNotIXDhoC2E7IW8RfA
uT8TM+7l7dPIqYWz5pTKbtjGLWSsvR9e63237rtDeqT5ibbUOZASYZoPvADTvDCq8D/NG41uNpDX
cef1Nqnh6cleFk3Sq7DKgmuroieYjWJO/TIlwlUW/akY9XDk4Tu3nEi+K3fzbHHImH+n5PGTRVCT
3Fyxj1L6U/z4DzOP7uwnGurbEALgDfjIfuT0zosa6+i6gt+YvPsoce8zbg8DhHSvveokO+oWfVBs
ZEpr3XCnxPFrqjyFjE7v4RkT+mLfv1zMskbzqSBi668XIZ9PoJWfeTZv6d9SxlHpXwWsVZaOyiDy
rJQTUD8bmtYuwjSHDktuP/zIa3SRjAYfPFuMEIN6aXCvl6WIqHGmHOH8E0JZijVsYEylMwVdUuTb
IiuR9Sn9ztXrQ9E8UQfVrZ6e8cWn/I9Q5EjtMryb7rwlQAOIJBdpA23nHCnCrdxOzqIOjYixiq8G
zVmke5lYY9tbGSztzB4FtRYTXwtD++sqNK/I9PDlyat4tU2n36XKKV6biEA+WznEXAXo68Q+BKNR
HZUd2FSZdLJeoI9OIoqyN45zJ2fri1/4Rg+U3ywRTs3iSxG0zVExsAkOWEVWBm8yGPCkTCmO6NVX
qar5rh5N+pxr8C+lfKq6/Zh56yxNCFsv1VA+Fd/u4hdVXcR9psDX2wRlmh32VtFPD3F8eUZg3HsM
afjyc7ExcDUNqR6We7BKsP2cq/ySleHofPHGYZYA9+uLMJnKHVK7C/tNMdK4YsJ7Qm+SIe/vZGtA
U3FHt6RgUbpB1zpVnxg6IFrHFHUEUjk6iLce2/YrfalNe6AbJV1KRb+wdB8ZGRrxnOpDAYZPj4Nn
U56JaToJczVVIUjGwMyNM/O6MPLulo7IivAYVxrkBKJhT8wwX8ELC6ZUdGfTvrjOSq6i8ksBIALe
bHmS4zh1bDwvJUKSuTDf+9cgieYhz7VIST2bj0NpNH4GYp7UPrqRS1eeaTIv3LQZnyY9aZ9EUbWh
Hhyj2/0Ee3SL1+SjgmRewilRQCEhT6hZ2VK8vu8rgpF12jMCaQvilsX2wdn4xwUnC/G0PIVk4cBO
HKDxQ1G7TX7H3LeeKZdzujLiEyLu90LF0V7DhxMlooD7OPL9r6z66j2oOFDBCVSaLzxBbmwtsjRv
2TMiZdPu+xgk2uQN6gJEXiMcNHWrQfKwoOXvs79eeXGPyfqKjJrK6i9e2LD0+AlfW4Reo1n5D3OE
1MrtCg/1rqQCsvquf2whmbBHBaEhv8FNBLfUr+SaYDhAmdPh0AmmqnfEyJECQ/UsLDnbYTsLRfaB
B1xdS8NgCvBa13P2Co6vPU+lrnNxMR4cVyiWffmbKWo3aW6t7kUbfUOXFT5b/OSztljIaxKKzVKl
+OyqkV6CIVKukcHOQIgs5Mq3S3grEJoLDDNOjKru2KNFaUfVz18oOofEZT4/QJ13lvd+bQJ20bIl
/rwr1Xms9aU1vu0OGsSd42vVNjfi5mBMKqfkf14hHbRlKTmtBvHTouQXBSodrci+rtLJ6nlCmvk8
uRO5YteITk3atPXcwjZ5ypqtC6/P3bV/yVa7ma2x9wYBB4uhWuShWQNWoofaf83PwBKeISb4HUQy
CVxrI5wKRtbDnPowELqWOYtEPlPcMlFaKVvKHVwoSNyZE9PGh29MhwGQck0VObapU3Ljn3sXTEcK
F7IkjuBwaVEc2Kq4xudfpUjJuiwjtzrbdKRoHs7nWRlonBItjnzIyWLplBuCdr7B7e64d/OowWy2
jiXzgdUZJAlSqoKe6SUrdNZEMNAFr+rxizJ8BTkDZ9mL9iuy5W+WZTQvAGs3+Ko/L9AwsoGhQV1o
UkHM83xia8ndOPrrOkyAQNDVveDt5TeKokJlaTw2VBafQgm/KDMfPgX9tzM6DBcZZeUAQPy3yA0v
Otnc+xOEtEov/TJ+HAfAaLE1+Y3l0arhoJVhOHiOd8OP4DFIqivHndYY0FUEC9CTwBMiBAAC3KUy
rWHiNegLPg6ASGodw8iBvjTSjr6uaxTfXwX9Y0KlwEIdCOFbyGiAYqdy6yzwbwULpDXxDh7BoZqX
sETP6rJF0em4uCdeav5pLYCJz9VgXzCcS1ud2fCRMgMz/tiHPK8Qt06w+Q7Xy3lY31n34Jyjo3s7
mWXNOSRFGi6XcikxaC0AURYuTCjbNBaIqKQSfyGrO6YXB5r0JLhoeM0sVCsepkIC7wcFU788Q075
ESxDrVopnswltpRb41ol67e/04TQOUeU1Apl/pY+bFlq3wCqOFZvfdX48WwI/cnbEsEvQK7vLXhN
yMGJErrlZyCVXxY11VGbNrLSqupwzM/fm9C+t6aDWs/YbGzu0oqa17DdmlmGIiJOyyPfJ3tiZmfv
ugUXCYvJh8fBfyLKY1omSLPLpCKyAWQP9fmA3giqO5fVnQ+0x1HkDdy8XzCdqzYRvtiC12YJ/XRu
OH1sBoNjGNEZ1cRqKwoY1bJGdOhzHUhCBK52vVJ9unyxfI4YijVXzKmuZaXmq2pE8o3P0MMu6lfR
GcIr+X8vYrQeG9SkJ1QV4XifhIhKfMSjBB6RWfyCd/YF7c+JkehepfPfrNRwZJqwl0MMTTMEGIQn
2LSJ4OXj9iA9WAVknRIw7KbDe1mAM+KZ4yIGqP+z39PzzuBsS/3iEqyKKOW8KajgkY0/5ay3ssdm
IP8j00qln1FWrswWQnavVkZN9MNza1FeNQdi5qP2VLI3f0bgINtzwRxMa1UxF530JZvR5KLxi1L3
d3ZFnj4Xrt9iEvVLCBViaaBlWuFaHu7SbzwPcoQcYlk9TqRbBW+eJLj+k/+J5x2bh7nhzZbEyOm7
J14ecj6oojRE/Kcli5X1dTatBo4xsJLeg5hL4aValSqJnqGx3TohGnbjtyzVuDevBQtg4NmARLFC
wzIdzYUVLfjN6uPW/G4+izpOPs33gOcyTZUq048kn3AxKrxylONiFngx+ZFZoUK7FlSQcHODefXA
75M7wUZvR6LPqWkzo44HE7mUOKVME7Hm84oOw+GOanwW1MePYigK5Z0QJTRpr7yLhqZLUXU5CVom
oI27yBdxZQrP2MJEaVsNgL6TL7SGJVB6RXDGikuX1CS2jz2+IJt6NGUuQsm22wad2McKCfmuAGVz
HMWPGZJe65rsaRzqf4Pop9BG/yUasphCTPEOjyr0rArN0LI8m3xMcfKh8C2KdrU75DlffMJSxmpA
m5UbpT7+b5dFcS0bMxS/sLHKBFyjGkXSPAZTAOR2S4iPb+b4UrXwGvVHizKk8bipY089XECa1mo4
pENWd5Rifk40KwXITtjKi8IQ6f7AQc38RaxdzArSemisiZBk2F7gvvsq+vHwKw03Ru0XxpyoVzXN
M0XnWdqdeGOswX0B6GENHL5uWmB5aZ5VDifFDrQOJBnsGWSfMHzQM95Q5EQ+5kiP961N6ZmnoV5q
+D9w+XVfwvEwjDnRs2BzgUgzG3OhjCcpLoW/B4zl4CAgMg2VeZIGVGOvY5dBhUUR6lY1zFYtCnTx
i6MnCRs9nC/J6McxtGOBF9CcY826VmNm5qRmtzBz3sfUe1P9P30EIUm/Nqwc6Ba23a6FUY0qm1OB
4k6e4UBM5KeqA96L6DdRIJ18AFFt1kVFIF8ejDWCwzSj+YJco5EXt16KfePtYmXi9joar77lwRMg
4t/dXxS/c4DBV8Z62vEHJVSgax6r0ln64bMEkwCgDsz/2CVKHv29PmArKhcqlIxijG5UaavhyrZp
oIs4okd+TDd6/lDlX/GQLGVeIVbYSWUQH/tAlc00RbuWR1JsuR8bJ+EkMdl0avRnVA7pC3kVbVei
9QIskwXMo5u4kmhJcfaPQJcAQ3CG00YKhTwqtQHOeuCgIL0aX9h0tlmmYstXldc8xEO4CL7ASv1k
0gOh0iyYPeahXEc6jhev5lffxbaDTOPKcfYU1UzPh9d1ZYqeHqa1D/ytCgJp2WtM++MDIg16OTJ8
MX/2flD//N99KlfG7T/7esGsSv+SUTNxaRClbakwSeERSIkwBhzLohqGR+9O6Xa/Vs8f2lqX2+wl
9ZnY3SVX/bNLFfFsZFcw6IGi+2xrsLfmxxTY4muk3vxFBRLTZwWJ00dBMf7PWTEAWdHc7sIFv/ds
1Dul5mkrY25TqcfItOFZCYrE9An1hAb56tXZ8QGCfb5tS8KmbSraGgoU5V7V4V/xfzyt8MofpAaD
4hGGCVuCREks9SM0OgJHrGWtBl6yTigJCoOfg8MVQme1BIqt8B5CXGZ5H5yInnpw81MXfnTLfzFp
7DbM79m0hNToMeJXMd5D9SoCL4xKCmSDX95IwZeaSbGvkPgNGmBe1oPCFE4R+OD1UxIIXihW1CTY
pn0SHbRVZ8ZfYOuu5kpyxcUg9t2EMtp7WEP9DcFvTFfjTCGjFy1DLVuqKFJoyBIOvDrlJSFC7a0W
7N7tcqVtBNTtEwWiGIYV9BdPgmR5V+OnPXi0wI56d2DGsPOmN4YUopwqAqRvhw4ZY7tmCw9959zr
FZLOvNOjGxhJcL2S/Vzx2lkdT9KnZAwyOWEXJ0duHdgTcfkGVt4AxNpXVr68WsxJf+uq0AwYRvkw
ORDusHKMy1LycG+q9pAFClWsUnEHukN39IsvTuK01/awUm2WPXyuDtqm7xZ7KFi4Z23XDJZAWgVS
8ptXhf0hGR6d7WU3crRtBuFqUMTYm1F57UxzTQghZLHYa9pV62aUG7VGqnQwkZ41WEOqEMLgfFha
W+BNPkIUsHPrSxFhCiIFctJ8/zh8qNuPqOOW46Zuu2xTK6aUM5V3c27o/6lVOj/oImLyYVTdVLLg
LGLsx6qiFEBBWu6JgSfNXkd8mLKs21M+ree7FZrlFDPeneHc3TA6CdqKneH+op9K1LeZ0o7Imhv1
dA0uTBw10lu2b5Cl3SSrEG80kCiiMWq8lsvZSeglfkYWkrMyA7cFhy5+Pu3i7urF617nygrXLJdk
yfwdNUk9GUBS/E+TipRGROxZppGsINZb2n+CG2bDNDsUQq2ymZ15wNvRXmZKfJMaC3YfUs1omzi/
XRtyMLNKYxN2Tz6V0l87Wpbhnb9HjqPyxMQzEtSGNUgcMKXpGqKN0QncqFgx4tyQSpafQbsqE41x
9HDemCmIk61LA5UXIJkZwXd+hV7ediSKaOk2tS7VjH7fo8TgSf5039Nft9l8fOhAraAG5ID4XjpF
T4symGedt3/L9xlVIfHwiaPtQyY2IZLQGWK92bFMnEczG7XW/XY9/tcikoJNizoFcR5sLL3hNQgp
VL/+beh/f66GwrS6iUxKpdYO0Nu95jZBqaP2ITCH6scoNEa/7KMEwDVH9Vm5NVNmCFRZJ1spWdiC
e4LBzEP5ftwhujPAMoV9AsAj5kkussUlQLWs1W1l12Zrvi8F2lALInHhY4ugA/pNCbGrBTKv4Xs+
mB3A8PCfuKedJt5I4mfldxqEDpw7imlazw2jJUDNYqpii8TokZycLkg8F1xmdwnpPaKA/iCV2dzW
gv87WpLLCoSilg+yO6eh164ZUDD74e4hQA9p5H8DQpDEpJLOTxyvn/NOj4Aoq5GTHzRRICA86dWq
rc0OOshqNbCBtbaWzfFmxj4KiPWK9XiydXUwsoRGLqrlz6HJxW1uLmI1os8q8Q/tTAOthDYJSy0t
HmMU34p0bbdOqfOiLj/Zv9rWlycvkG5cQjYqBX9C0Fqhkfy0u7ja52FpK2YRIwwKrpBkxaERjWU9
8dl97pHjHysqGMIVqK6wTBKVUB1IsEvCEX1Wx+snyZ6q+zrEbWXAo9Lrqnp4deQFAdK7OQnpHzq6
OFuWMGwIXV2NXATnwGwGnZJ5m9TlWZC4u3pN0VFaJUUfRVDdiKVjVrt42vutxyDh+L/lGPT9zj2c
ZWEst412O6nUmKjo+NTEPOIKMr8eD0qfjZfvQH66A71Y2Xa1GRViPjn/L5TDbN0GAWpThoZEjlEB
SKkGlBEeSNaXSVZ2OjPcVxXd1jC/xSMNUVwR1FfRcGF8xo3YKbEfMoJs46KWojfGo1BTcJiA6EWj
OYUIgoH5LUXkB5fJib3np3AFoawFlLf4tqYoC9+sFDvnFx0+SN34Tv2mL0R0sS0UuKEvXr1Jhd7A
GM2vEdLGM7wPTwmr8O+m85mS3/39i92fgXsMwkWJmoxaSH2hRgpp1Xpmxb1fgxfd9T2YnPoaYPWw
f4wZSDPqzt048jm/tRnwtT9lIwZnvAvlBvT7s2H459ke3LYZIz4LcEw+ZQSKgpreT90xQH6X1fwg
iMVI8shtHN4O707QHCKsLaLYXetCMkT/1fnmrexPzCyOfFOU+6ZbExgTAlGtu4FoZjame8tA2bCK
nuXixP07xNbtYfDlYNJASNpCCwxpiUoGs1Otl7zozSJaErkCXjSRf4ABhOT812bcXXWdwZZYaeNo
1wDz1BJD+1XjgnqHeIeOyom0Ak69INQeLbWPuj0mfmZ+e9zpQeTYYy4oPfQxoEmxfgxpfUJF7Pg5
Jvn2ATLvcg6ej82EcTL8MbVOjDm2U60q1fZzsGnQCPA2VySJy9r/nTHef7zhjHRpH7C6R/EIFczx
L5npl/2jNGWWBUI0NDbWhKBQhzBaNkhTcv6eVSeh3JRv4o8ko3AUGE3Hv0azp9N51n4I4o9XICpn
lkr97Ms2QUxbyjtJJB+oWPM2GZFO3ag98l2vS/efrTIj4+4UV/la8flefA1LTbde4yfSMwUUSPcd
onT83KMzF+C/ap2R9veHK0l+Z9d1BsbE09Hywex72grpTVMiA8LgziNxIeRUYUzclyEarna+Fipe
jG1BBxqb5Q9O7I3/Gq0uElSc1Po5UbN4AEOaZ7lA+q0X1OPWwKXJs6dprS+PslVasIM23/7xGqNX
CMmJoRG7FaABp9Ie7ydlQ9CdLmVwEdLlH8NHWvcVIgqtYZ4JIC0YrReUNrEKCEnqm+ClnhdTEPgu
AYV5OfZi0B6vuUPCtmIfR09Ox32aaIKW7qQx7beTxLeDKEiKrf/vwvYGTvLvaf/YgWXXmGMV5NkK
3Jbjz23VQ+/MHir/4B6Kr1lk5T3A3C9xFAkkfGXNpRGTRP93aiT14nPAYplqOmfyhewXn+nP4D8y
mjcwPhGWUt+53+Fi1iFgjqWRfg16CizW0USWhjpxdbpAqH4zBZQH2EN8Sim16rWJGB8lQC7b0XwW
QJicNt2jnyd0CNks9AenaMUgKse4wbeFfONQQncJOsUosGem941ScKWRlexbirdEa7Qcoonsfij2
7j7/BymWMP9YyV28xQAd1lfo8ERYhB+Cc8YX8n7O5n+Uv8bRAV0CAkjUJVhf3C/xfFgsqxj+kwuD
5OnJgoLxw1VUPX4x2SIxUwbVGLQFvJKeUJ06Y4lwlNBehar94hkJ1Jbfl5xOGAGpkr47Wx3vcqRY
FCe5udXMPfyjW/i47CdI2A17FPqws+KNg2pFXHU2dGIt1ThfRYt1/nSL5u+0t2DaNHzdfTt5mU7m
DZINB3bqNHPpclP3wZYATl7wAhy9QF9DZY8fmlQiblNrLttlKhpux9EOuBg2nsM9gYiQRTpxdJcR
TkiZPAbIAGvounA4KX4C0yvB2h0jc3xZR3fTIvi2Ngxj1dnbOdkd2D4sqjjdPZgt0NCXFBx8a/be
xDOW5NgdltJoS2Iiu2Iod7qwfE/mujt6WRUvvifhQLY7jGHTRMs26CI/kFWKa483Ol0qoEbEtUbb
fiAxKl38OfprB1gbcEOhXwst2WDnLSaG1zYXMzPoshDzSJiETj4Yd7zAj/zZYYCYOwIu58mcGqxH
v3C+O0H5Zn3HCGz10ghejMvgeIKmfg3eOn7pX/qsuTc3nChokzg3My9p584ZGVIW307/fn1mOXtI
LdRDpNme9x7RhnFHMJbfw1egURxaAnozOeLXlLaLtdLSOO8bCY2pWffD3td2a/mThMfcV0wzRBV+
0IxjRRcQATq9x/NLeb8off79Q/goDoLIRqOsQlWOYhE2jcqDvZdCxq1/+ih2CMdhOGsTGw+fLJEI
jSPe54ST3oBL78P/Mj0bBLiBtN7Sc6AubdwcFLMH5RrO76fcDEi4RjZo7NP9NF2e0T0C25zMc3R6
OFbMircNZZ8A9RnewZozKvK6x6sMfjvgumKYKW7xQY8reaJpdicrkPvGyV1kw8rSo8+EQ5PCDoaZ
COredFPwYrkT1AzYr+76M17NnGgb5Pj1u5tRUxIsoy8kVQ5aCS9rFiyWrxyiTYRCQliiP/Zyysob
heyHuB1P/6aZcc9Dpr/MDOz7RtA4t5G2VLe2QP3fa8+QY6hwMcMqDMlq2U1DNtG5VEomoxTp+JCY
uOJEHn5QvyyF7zfaWM9FqigqN6Fhe2p0oaLFoGA1mrvof/g9aUS2DYGVWkVrs5W6AV+f+MBb4Uww
M//eGkYKuRTbTUrM3Sp8UUDkiZ3D3MVA2Lyo6tKhDbe5fe9IivNYFqiygTTnywmK+kj003vVkGam
b8lh+SRIpxRCmpXHayhhU1NjICEv5I6E6D2rQfsIFMoZJyW9Ijf1VgJNLkKUR8rKBvR+43exDvxy
HULXp4o8ar2lgCsjgC1XwuUBNJ1+A/yrZ8sV6EoWaOiweA56DK79kShHHvDtUZbo2ryxWg3btItb
11DWTBGEHPr45qJW6zJdanvrMtlZsRM19Quh++kuAOp9QbXSPRMva+CCT0DHqBe9PNMAObLNG1Rj
Z/mE5hr0wYVj9li5kLt9UGtNZ7hR/p51AjD8cakH0TmRacR7YD1vnnRpKn7Yra5eXGE+D5QCKLPw
v3ecblbuDRDQQPtlkZtUNU7n8uKv+pwDaVzurMMtWFfPLpLUOtlnR7AKFZkwQER7XfMFhgkQAGyw
6+tWwkpCjdMbYt+/Ux9tQt+wk6fAJVc4X0kZgkFLlz3dvA8hJpHX4rtRo3VxyfGlw3hwRZvW+O3O
K8VveEdBwZIWw1w7cAOetdqurz6nauLmZnXPT8xocgKyKkwsfwBOmBgC6V2SDdQYBmOR9Gsk+k/5
uGNncKusvKLCjE/LB/5AdqH+wwu2uoODPyidJL/vmmaxxVX6wTx6cab6Ah0AeIydJ+++ptpLObXm
SeR8dfEaz04lM+JG34ZeFoGnKqoLM/RK3kvU8bpr7CmYPFh/FkMFQAG8HFGi4PDtUhn5XyfvDMep
Fw9XPFY7vipGQ467adFrckjIpod0RX+3t61rrd23F07Fj9k/kw/f8ZnNrO4ayXY0nJNOXhW5NVUM
9Y7gx7JleFt+8MYkXiTryK+Gxs9huPDBlHnmXTckmmggkzPtSdY84vaIOekLKdK+e0UCpXasNMoH
qc9KjnDfKHi6+0b9QcwZGfoDoF+mKrtmPgapgdhe4E+uEYwrWlz5QbPM28tOAvKO7i/dtA1zbKBd
eeIyLjPDQtEc+RJTAWttFRE9jyxkrW7IIZlkcHti9+eVzsAbopvCDxcH+N5D7N9xwfxNJ16JMcKa
ILI/azJQ6Gz/3oTiOna8scGW2bmyOUiUHYsfs+QiNi9QgnChTgNBdMzRpEvIOOvHXoaTpw2dsn1J
jr6IQ4PjxQnIVMAuJ0MN64c1Ae+RB5smKsf7c8PLSc+Nz1UpW2ngo5nTtpok2SUMRMc71ZP5Wobw
no/x/G0eGN9hgTymI3H31Aahk7akzQNsNslYN/O1LqAANoTBN/yujh0DRn8sawC4Tjfp+VR8ztOM
VmtawOB/MevJv0t3HIs3PWRksnQEA99FQgx86O91xguCGWFcjWaPXIdum53OWravbjcGO8CyfXel
n1a3PUDh8ZicRbWUDJroyHXP3nxUrBdpvOs/7B6Tr8WLHe8rV/GO+4qz2d3CFsv2JOpYTezSyuRS
xep3AUu5M51ePnMZlWIaXLcqW4E37sfsA+zzcRdLbJd6pZgNo7d2yxesV/pvkNwwhU0NP/ZWbjfC
ro20wgDDu26FzNubMmhI2vCIJH/j+BwX0FK5WP3NFcxInQuYgTz0vlG6+Lfo9FjA5AZWfXlkr5bS
v/79/Yl+OmMM3MiSMjGKsI/2kG2BA/8M6sQDqekV1Xq4151nQN7Rx1dGyvwbN/CyC3PJketipDdA
qfMZBsIcBy/yGroYr8RsmxDZdS5J4wXR9V2K89Gtk3Ko6eeq9xJIHwbxz8clLW/YGhMSLOD7Yhm8
e4pu71KvWe/HoXeilNHW9o6/gq3l14gHzInmxMMQyX+sCTjZLZjzpNs2OnWM/h7RysGFIu+qpqkU
3F4v6AuVacdjkvXOv/0Yxh94o+9zW/gdO9YshQN1J51IliQvZK9Vwm+KcIEjiO84PiwzVDBJ1uTX
if++wdDLU1G31zyJ9spA93zzEHHXr8NRJYz2yNp4Smxo9+VpDSFuHnQCX2gujQ5lrLiggFMjDJ6S
/h9geM7bM8xfZMxX1F7rSpnsxI6E7KQU12J1gIJAFbBhZptcD0pzmLgSift/vl0cd3gvXuckq7YU
Wlz7rzFAI7GZAvtY6P1/F9HDMFwe2TbH2vLoFNdzDqRnBn51E6++bD276zp806HYpBAGHQNuP5mK
lHHJjzX5YR/jqJOmGsLYRIgDjxZrkzWeqJfHvV8ZEb5wQdVHv7amjgX2bSTJe+ZmWirH1xGa7K3U
6Aj2B85POc+iO9+sx+EdO+3LJvcn77tb45tMgCthyI5DKSH9OB4n/bk+5UyqmaHOo7TGE+2ZtB3N
/fx9Ppe5jojgd1Ys7MRRaptQ+o++M6u7Eg9zQ/XRD0KOdod2CUkotlOT/6leIw7GktMUEQJOHQvb
DQ9Lbbw9BEjJOYluT0GPZB8HdwirgFJicFID7Z434p0mwQ+XCOcPy4tt3156BBca7pUDUT+ZNE1D
0q0ccLXaKTWXXUdcXCuuj1qXKvMKsX3YTendlUI1FtpreIrBxZjbC6XLMFl2a7VfAoR4oBJqbYrp
g/wgKUIrP8yKmlrlcgpVHq04CA4/T9VMidp482edy22lmH3RsYhraKFjUtcRT4RBuUWGs5bJ7F3M
sT2P08T58uom/uiJ+gwTTUReX/JFNeyutOB+uRd/RjAYwMCAuvc/oHVLw/XwDAgJXY2UBUK2dK4l
rjE48TcnNQzqWRNDUnkz0H9ugl8j5ne6VILGyQrxACgFz85mYqvg7Tz1HqRuYB5geBlXxDsjRqUD
BbHSiLSJfUrewxYldpv6QnmFn+utBFAHqf40jbcXyUjy36QfWW4/ThnO2SpFHIp7m6DC9lf+xsbP
GaH9BNTRRrYoMi1GbZ/Nv9lpEHb575eMaF/SWs0ghevfN1leoHB55MmwRH6UnriE5UkhoGFDuLWa
1mNdNZx4Fodc1Ydr77LtC3BnYmgUYmQSrpikKUW/Gv7Zi8+cZe3yU4FcyRHsBcCq6hiVmKw+5jCP
Ao1laUXsukuk8jGiAW4rYTf3IPRfR4mRHpVf7EhUglai6JWzdiiWE/IaoY3hSmx1JigiOKlA3Sa+
BLUbtEkowyXJBa+ZqPzMxlRABH9IY5ErsbTk4c2SwMS15yONyrpK4r2Y5mHcUAFH61TpW7Ng+54K
pageD4xcxX7UWoZ1kmn33wAsDk6z65P9rqZOwfIIn0XynHjKCYH5Y/8CorJ9IfthyFzihEqtF5LF
cnwjmNf6hyQ7eENHT58t7xzIkKD2TL3knIOiTVnEqtsqM3prZ4giukwJ4dBJwFb0Bp5uxoAo6Q9g
QeCmWD7V2WEzf3iW78svvbHrkg6iufFX8wSR+FRi8+w7x6x/4PtQT4HNQAQKQH9ucwbz1aH2uBgD
Ki7LgVGS5jz4Hp17T5ia4ze2UVikNAHRZnUHbI6Ll9mN/n3uIYKxjVrFS/7bZ7iUrYJzveWEz29e
bWVqOxYDm5z5lGZSFbfEI88GQsbyBEoK2BYXEv2cA617dXWvsrKfWEj/MuMkgD8wgmeBbua3sQoO
+SNeXUFta3X8JIK+xvcoaq9W+jq43+ysiisUTyV6YIzISdoS3BI4f5cFn5/gLAqrbPsd2urkFyou
KG9SRylR3YiVwkulo5tBIKZDMDP7VK7I+r3t/m8oAPHWUr8IwOT7Dz0+LEsaKYd+zGL+2FXby/ec
d6A8ccUbFlVp8uscOHbgfX9EKYMhgXRDjj/EdMwLalshJJNwppRJpnRN4Ds2+mb995+rPysBUgTa
p056MrB736j90EpkWqtnN9r12/M+l4AV3fqFvTInWWWGs//KtWgVkMvLHj5w8ATPVWKl08Un3+b7
hoyyeZMc4DLe8uKGHpr1cOOL1n2LUP++TXxFdjs4UrFI1dTIm/UtN4NdzoqLzKVHqITUJS7cTuut
IyhF08VRhvoxgf77c1jXaXpC1tVy+1QmMDPOlYybqDQAk27FnFCLsRhwBQadu8JrAD285ie+EDoe
kO6vVs8yZZZ/EG0dbydDtbDSf3oLHY+tqMV58/Txj3mhLJG8X+WOSHakQHCVafwHZTjGomdNE0cN
w7g0mUpxkf1k5WB/e0Tf6Sg4NfoEsru+w/JDFsv5RbNRs3GoqM1smpMJ8js9LUWU1FAUCiK6EMEx
5Ty/RCqbKp5UUOJveqjxjbuCw6lxH4GPcV/eYcRmIH/VzqTd+xgZ4Gi7C8npwzexuUCzICzQdKWB
JrpVB9UbEuzBsYZVVzPNAmdT1phGuiqBOTTBR3chAAkfQd51CkJaIaXCM8+fNNfMtkUL7Yc/Mf4G
dXwvcSg+sOEEerMpPOv3lRh7peMl7Qo+WWX6Vt0SfsT89QKfgvGkoR51FQNXQtVf8pc7pWhET5ye
+TqFpHFCV33MmoNSkumscgrs9amSDFvVw2HJQTNZSoJb2JiWXnLooe7DqB+nRP5XGKFINfwlrfUI
d/yo/0wAK/YJRBj7lyZuY2KwKHiIRuHeh0H98a6I5sxc7m1/J5wutsQ7rBLQUDOYB9NGHLa/K8eV
NA50O8px5Z/d3iis3cymg0FXOoWs4qX96MS2AqjGv2iXqRvJ99VdirxBESpSKRYrJnU2R6eDcwyl
xg6BTuVKmj8wwToH6ws8EMCqrsA0+oxQu4pPP4qbEKoW/+OLbXriBH9H1Lc2GQsUMaMYJPlzMWna
G2MAc/f6CyeaLUjr7CJ/j1wF84byovdbat9N4Pw01kY98WTn+wR6zOSZMKUQE+N9MvKu4gPNwiYf
MDbAmxBe6MsCqthyjKbaL0n1SGb0rSxqkxuqkbuOvn3oTjv4JTrZknXItI056REI5HuMneQpMUgs
ZmPyQH1F1EQ4MB2efuTJViK5NH7SFXZrcdKSwTp2kjlTw3ffZEPAesTVq+CNWZsfwnUjb0NfZY1F
DSR9gPnjE4p2X8oJT7U5PKLSyZvdN1xNA3qyiX1ltGs8wn6rUgX8Ot316tiY3JWiCmx8RZjarWRw
U8qNWSMFlFbJeq10lkhlHLuMd/bvxKMFudJbocp2r7fwcwdJ+W2ZPqaOHQiCi63nIYpLWa2ZDdv7
WcgrmrQ4BjZa26+Q0IxByG1iWCZDXBblF/vndejOZ3RU4WROVL6YGXRQSilx1O9jRY7IOW677cCl
Kec9xqtnNvXPYQOFJS+1S1Wd4zJ8k1L9cF7snw2eR0pOdic8sen3S6JYQ1E857G4ORGq1V8B97/c
MUs55WwtPclFah6AvVE7rS0+Kd0UBTZ4XPaccgmyOKAsO1Zdyhu2GC9p7ZurhaiHft9lHlI6nB9G
NvxKU/jifsiS2RA1soOzRcS+SlrkCc73Yyc4aaVA9ZXZL1nVORqmfpvpzQkt0bYG5Rm5JmZWEWX+
DaZLn1G2syb3MWEzxsRtsGNxWZEFp/A7MVM4lHDf4MSXdRj+p0jcZ6qsn8Vez8Xoz7aQfOV3q8HX
H4+jeCUMdOvyZFidAJrYqmrg6bqlLxQQE0rdNVQOqdMo5sqS5QLVsgkIrs92QIRs9z0RRcUpFIb9
2F63BskKf03N0CpEimee/ZDUI4MJeuKHrZLVg8Cea98vwLp+LgA7gdAsYLusxv7ANr5wo7K3VH7d
z/4U2Ntny8LNl+SksNBp4v0jnZeggMtyUeWNZxQpMC/i6k5Z0EYbRPk5c6T87PcZedk1c6V0fmv6
x4fo9tlt6365XoDV/xPC4XGf5jJFztksZv9s8LUzmXeGpNjTBTdQ8EB2uSp/zz4mluOzm34Xjwu/
hGrg+rby92PN8aqa7G4ciOSxkd6oCe4llgZbJ0nuHIcvIWTk6r05dKYpqvS81yaQb8nRQl0sRcu7
5fSHgBsVLcS7sbamz0TXisXimW5dn7wTF0KWB/Xa/ikBKdxLBo3ic14y2XdtkYAhEDt7zB1QE5CW
TIBnls7LzUkAtCtcpNlnvoH+rpUCR/L9elj7ogwkrY1EJWhXtOCcMMA/q7omOZ5wtM83TDYdfXLV
ddu4M0VU++aNbAzuPSVTfLgXnOaD+CTWz49ndpiMGyxf9y3iIDvU5BgPFWaf/n2cHSMi5juvLZJu
3a90zP90LHh9o9ktmPEQsV4cW4W3Rrxk1qINL6L3bMIk4EBkGCSLhrGwRNX5YR5t2gLEjkWkkdoH
7N9oA9Zvrb3t77bHJxRrur+XoSwKd5P4Lmd+xkjAEC1yeZsKdiJbIXJ57IQMVLun+6tNn/VJFwDd
4btrNKfM2BdcH6IIKLfPQXzyc/q1Bqyq5TlJXKkKWFUk9wdnHShUSpdqQd3DwwlHcRabuUsBRJ5/
SvAEpb4pjAlHwNIaseNtns3rwUferRJ99qk6s9/I9Pky5/PeZ1Q31JJ29wZ/oir/N5A05iQSGl1U
FW0nAlA2IcVgZy273V7PePlwIohjJlWJ9dcmGTqdJlLBer/OOlMb+fifEfPWvgZnkVVKbrfMW1lv
XShITwKUfxe9c4KVbzzW9a3JsyV3Z20uWDCyq4SHRlkK2Frp3TRjvrsk02UKXD2NQXCNTL2eIdT4
m3wDHdPc/LA5CYJJo7zyL3K/qUXTvpyStC8nRlH9M+sAkdoju6OvVUs+sPUDYoVcCjaVjgEnoERw
sKt7o/sTX1WLSuw1NQKXZxFON4LegzzTcHIJF7EJW1gWFKGVhC63KGapw4x0GwfeWIUS4CFiylft
CDkZP+WpQJFVHupsyGBqFJCHs+Yl7x9YMzxJcUFpoqWuNgpvYkUse5Eyo8C5wo+c35Kw84HNyUMU
wzLJT7DqrT0JN9ufX+4hH4sZrCSFyLgRqoqYrW0lsvDrt7KUOrANgB5bcWxXjXxYjfF17LbPJ6Qp
mK+FH7OE+jfMQ1YREeaVzZstmEMccpwbWQqOFt7RUxT+FC0OQxOCnigPTtkPS350XDTqvlxDeSh5
bVKqTwJR1PNYN62j4BukrzHMrfT1XXprTwkMOv4bhcoRCv/uw6LUkmsh7Wx2RrUvGs8Eqs/yNoIk
U79ug8UCAZ3h1B+OyKtOW25iZjY96RlkY9dJJXU0iJwN3d1aKKMmO6u9FlBMdepsVaTozZnRIa4u
txIC3kMVjHfxXLFw7VlkOiQqURecJFnieokM5KdQEU+ZYZAKWVcBZ6nCXgwJQRMh/eP9POjnO3PF
lckuh12QJ9jymXkobV2xu98KlLGxOuNVCYrjuV82TEeOd2NC1Vl/lwkMaOM48EWJI4YlucG0mSrj
QDfDsgXNd7VI8kWfK6Elb+KLYv3gdOtunB6aVtjQkQxotwvrRcRZGC+Ek4dAcEkpOnk8BSwjkt7m
ZEsxR7MFS4CqJNZbOHCzwpaE1tk71RCIpFB5ryP4q9O58Ye+mw+syG+GtGVVoNx5V9oUFBaUBz+u
dH5L2AjF+lqWMwy5UOt8s/g+9IKOWQqj7WApL1Kk5Gu8/ruNY44QYAvkd5Pss0KnB6uCLEX6UrrV
PX6qTalls5HDG6fcC4CLzsGXsdL/zRI1Qgvnr3qk+palp715kF9ZBuQ3kPU2vR2dPO5hlLGm03tt
l6nO/G1NusMaCVlQ/yufQsnnhIhLvReZm6syDxgUoXf9pT6gwvQnBKaWBP0ibuPYOPghZZiqxaQT
cr9chW9fvXe8AOOhRtSGmnCprIX+RmKm8+JhPSrvrJoyL4+UoJX36lducJ3BMppP9hH/eEuMtSZg
3nPSffTxnk41WCBewA3Dk3x8Bnr0LAnmlVkMhRe6k6AEcOevY1l4FG+4DxjeCY3h2q0iFZ/GDx6r
NPhfcB9bWSRrUlZuBXO3qZEaVpnB1GD2w2iJCQpotVbGfoGTu6aY6PuiPzR6jEgql7/GXZU6WU3d
ADcYMKZKzV9+yZTYTppMLZUPPtzstOwDQi92f0i24Krdz5W1o4ktXy2LYfUZ5NNTSKfZwXxS+QxA
KzXMjBveEaV/Hp2uU0GvCByLez2On4KHAULAmKa661+gJes9/abdaqaTfc2FvFGGjLQ8LK0dwHNp
pLyBq/IbpFzI08i92zcxTichsAOrRysJ+IlG7awb07/Fj3lqY0armnXNWdw06kl4tandDZMu23Io
/BWIG88LzlJ7MlrGL43QQonAx0SpOmhnU07F/Wwk5gM3n7KTfXlltJRMqhmpNVS/48tQJKNS5HE1
oshWL26rHHOwpp3z8gwvPiPostBlBFEJ0n6QO3jRHZIAhS/d4XPpLJAg6ibPCeZdAw4zZZdNljnL
OgwmYK6ncDIMVlZMs5xrpXI0IQtb4bY/FNc+IQm8pw/ZOSXHhnq2lwTUw4/mAnRNnjrfTpHpgvNK
ZpFn8kvb9YkaXOjoevKDrXZVJ0ZGC3kM3wIx1IXTUr+fPQ76PjzL7NIjJR1y7DCYw5GUmZ3tyTmZ
i5QAjuM63Tm0eUs6SSCH8ryEVJupGAiY/Wyf9d/FBieLDkKg/fNmjiNpS8bvTjq/8qfYElNme31H
+QvZWLnnndKLm+4LO9xexaCacWA1yqUy16Jfse+BHarPqfoUcCuTcFYgdcmuCVKzWlLxlP4R4UGm
pGj+B+ugo1okIWlq/BfMazMPjh9ba+E0TxXMuwVzTDV+1dJYJTK3A/THp2XOZM+5Ip5tEaJljaaO
vehPAak2ysPu8lT+odVRhkYgvzGP+yVPgvkS7M2BYZiL8oc3hZiYaaaUHVHf/I8PumfKDDBPypc0
/KLrR2GpcNx6plkP1HerLN7F37U2sI0BprQRCc2su0TlhKahI29PaP4C6jDV7YtfrMh3xop8mFOy
nIHJzs53eg7zVVjQmnqd+huK5g/GrIxTlZlXfsTh82cPOdfy80d60gLh9YEHx7uIPmFvbg1kaTeT
M5Yl4mgyiCVrhlrgIBl5PnVKnQkFVIURbw+5yveeAebwxmcMOey+VEplz0J2y2ah6TAM9r29sfDT
yUpwL+PO12nwXbUBGJn8c5m4PqlI9j7VAKKk7ZTtXjTci/FzX9HoW1WfWPm7mIC5BHYsRUTEsQQ7
bLNDWW1IzhkUWLUD+F/jZ7aeSH5mx5NMjdLuBtpwCxjbUVZ8uxejsqCBm85Y8m39grIa+8SfuDP5
CHySNPDRv0Bg2eG1WfvzaJlSwDPf+EJtNUFGjKQIhzv228Xl818PPT8PKzS01HAPfBlQZFtQGxZc
KnLk3asla3lsQ8lIHPdqxBz7xTsrJJe1sQ/FcVX+afysrSQdMZn8F+Odu3A4HJUY4hgZw+j2Zxg/
7nwgDGqGGTKLP93Hl4X4rTSis3A/pW1Uz7Bc30VzBWrVWV/lf/P4XbKLsPN02UwW+jPCrzmgPgMY
RfWfG0qnmB+h+q0uv0KdimdYthtADZf4mekQ2G+BqVLZZakN1oY65/pJUGFeExPb1nEvwSr9r2U2
IRtAzxcIvI4zJa929WABHb2as69SN3o/LHz8WFjbZSSk01YSHYghqdlBvYa1ZTHCLJxCVhXPUCBD
WYK5Jku3AhTAy2E102asrkDUzCK611EuKmvuB5FX0tsMbkhdFgNSG9GtsjKuEe56pDlUkIXuB2HU
YjmyLthEo62krN3Ujn8kSktXJ6fs3p8X5+w5xkgfiOtuheolPNTTuvaXDSNbAuVuNzS3LfU2qr8p
T5n+LZ5DcG10xf6xoBkwkBJ+7qXx1joMYojG6dv5Wf8GfJ7Aid8CTMDVTEc+JAxD375v0zoNcppP
4FQ3W432PZhSrUPE2/SS3a4OqBQRgkFLNR1gzex9DTjfbTu6dxEn+e/ebX1c+KRglUxT3YhuIl7m
3HU/k+9JvLsVKgzsn31kgjQf8gKH9nVg8U6/WeqC+54xLLGOzPEkgxJTIvAysUD/wj3oNL1i+PM9
dmG6XUuK2qMA65O0twG04Et9O3a+OWOemSkEisX/y+cqWTcbnjwEQadhsPAibge4caqzgVCgKAGi
9D2+pRoDH21qhhy+HllbDn/sjfaDN8bOVuRTmrtNEjIne7jcbrmmb8P75QK5CuEJf17yMP0H9Eyh
puiVh0GScfSJupuWMKNo6YAxILtbVwXCoZ3oOPBTE0G8wJLtKRyc+WtXUJ4JShPzYLm+Tb/1vm0M
Ghw19ecS2fCPCxTn6TlQR0bf7kxRXrVT9cK9PSuDcqqv2EU9/eZaW8uaG8xmBzDqUHlL8Ov4/u6k
UBz4KFKc3K3v6WAKvfchwLqqbhx3ukgQOOt2tAcEaMcoqWKuSD1tbXFSnRaH2na/T9MoUSmRILrI
91Im1K3RnSo0OzhrhuS+8UD9PSotawhMRfKlvoi+zOkl9oXoJgfZKZr0Xnk9BJ4pcBpUbuo91oGH
BQfnFejC0eKIbfljHZyohcom5+/7qOaUmdehAeuu/AqA54UUZLNgvtdC9UTzl8ycaNeOtTfkZf0p
a6I8xYgNXoRku3yYKi3Op0E89L3CTOEnZOG590HqXawM2i4YjWNDST5TCPIWiVjgc3urFauRdYD2
aOI8qa2Lxctpg9ue2IoCl9/U5/JhMPFh0hQ1LTw/qeEAA2z02h9A+QVujWEV8xUXj6v9ORmHpzl7
DeAluOyRi5+3UjUJBdWZFHCMXg8UixHAN+bvEEKlcS9CkoDE9IqC8/sKcIhvYgb8PPVvBuuqgaRs
LiFqMp6Wl7BB/UnCgVDG8ap6EPfsfMcDiobkgirb3TyrwFLPQfhevUVNLzArwCskDiL0ACw39MV/
dzay61wh08Ww47ytWRXbrj/niau4MeD6vpbcFmcMh6YGCDoU7IrXQRgO/fyt0XTdDzmg52/Ds05u
mO0MlteA175fsIZIYMr4kp8Mau4I23NF61FyYQEXoSosJEROVwNpBMjg2DZPuCR0wSpDZCBeXukd
Q9iPEUl0YZGiZMXHun8cfe7kbvnXbWcK09VLKcGoMELFYkGc/Y3MWw3GPOrOyK9WA4MVboLxeiAF
cMy52YMd0sJ+u12km4Ta2S0zlJFJPUzQnNwtSuauCasNFr1gUGR3BjHbIt/aq9UJwnCLiWfwTs5T
FpHmfW/ovCsTT82/v1NBGSul578l6DJb4t5r4ER/Nj/VDPeVrzDjyDI0G9JilTgy/VMAV1jnVfoy
ZLOQs+z/sBIw6cDN1kMRBbkrH9q/TxDIKTju+Pq8OR+g+AdtQaIge93G11pnF1cIGH/OItvBvMWw
Vzv0Ayx70ZTtgaLPfDQqwx45sLFnZ2IVJL7zKnLPqP8qi78eEjkOY3ndr4UFsstmdVXWn1CRJ85n
IRpVRxD1FR1EFNRqgLorGef47ZtltICbte1XHVqRPDG1LlF8Qh/YR2KcLBvUUWy5XDfuAUGOr/b5
2aihWbUpZmw4mHfJoKcuY/3lPj8jmmXC+6cajEIAud7E1zcwTbH/WR57ZrV5QOMNCzmYJspyE1Ul
UuibP2H3+iA/Z32WJafUsu1KHKr1PZ9Hn04WT8U0Jg7ZTMmoUrbxT4tAiCSzzvqI3qrcIGC74Mqc
xOg+kxvtwljF7Fe41sujUKmCtuPrkFbW6spx6BZZraN9qqfAmI9zeeFdaOluAPYZzB4qUVQdTMUG
pFgykQdRcBCQkhF9FijWZlPA1s37x8/zlZQECtgYhjNwdNwro/pn8vfI2Lp7RqbMrZxHIAHYMnN5
9yFx+MvDL8JCkIrpP8q1PBst4+hBZbD015uyUc/2K6Oc7kZQJaY5Zlr9jCTC/P778xH2ExW+sdox
ZacsXgObBPqq/9Tv+bilaiL58np1h5ECPovaejbHORSD8Dq6p/rkMSjfMidPTpeh9JYX7TuBknkz
m/QCp6ljarYzwrIe7yUiWQP5+S1vaZ64DH5hRsoSjrsOK7zocaeLxUjI/XFLCJ125BB1RESnoXao
Og+28PY+ersdjcmzNZiFoQWE9/uaJy/5ToI7CPNbaSYchofAsETAkyewXm/paw97dQ8heqfEO19b
a4bTH2hm9dJBej1U4hWHQ7VJEp6yMNXJRdLSJ0AQnctN2ml1C5RwRcAMMW0Wu/fCRgcfNVm+NiDC
tfIDDJn33OEl77w++6UyjV99HscRvfAelOda92oPxgbZy4N3tw9EhIhJp0laVpKLhiZvLW2YpkW2
9Cqg1Ay+zvfLwRIlpO+ux756aiu63eCCLrfYOoDR3FK3zULiz69efPrFc+iSfTAMzBatfN0ti7iH
aInIGrBaPcj89dn4FDJkR4fqe04CKIhFTkwEiu888dcAOhFjNQvwGj7YFXy1ZcFtv7REEvPTtAvN
oTgh8DAE96z2KwDPBxGadGf6GwDKqYgy1M4QPIP1KMO82L5aYf0bnQrHP0LgiBQl4SuvFurQ2TD9
bnNLRcGpmzEb9535VpwHueduVjNmemWjg0PNTbLzEwH8tYHcZkTpoHZsEiA/jy/qG9gcnPDkWg8v
kokxI9QO3y2rzZcErd0c5jd42yYwK8ZjR/4xxYdlFJJy4YP3L1ZkkKMyI2bAMMivOFR6ZFH7T0rs
A56AqmGhpaKj0gjem9WYA4SXo5wNanV53eIoRbeMEHawWhAHNo8xVUJ4MlnJwiQVwwgh+3MJiZOU
Pwe0QS18U4JFNR8ZY/jsjPqMLhd4J5sjR9rSTLzDlfDs7W9pDGnjB4jliNZAU+zHzZMUGByFGMj2
m6lV0XlmGIXCy7UdoAHz2qMaeHOyIkyNFVTzmubhK7lhm26iRhTAZVVd0RIkAXAenqMEttOH6wm0
5p61eV5cCAIOMz+UsLV9PUYBKvYPBSIrtTNnL3CwX2fBPdO+yN6hMx0iiVO7p4L6oiolkFPy6uX5
1er9TBjbOSnguBsO83mQx3PMbFxHpNcYOa5gGy2WfaIDXp6AmyO/zn9MnoL9b8ks40fjjOEMKPA8
A+wdjDNZzaABQxpNOIePghkEvU3iF8CJfnCna0PxthU9Zi5fw59I8ptBAQhsxXdEJBg9uUvZIp6a
cURHxicwGxjrceHj7VH0LgdTDUAwhqBGXBYRLq8698BdyAT+MFsx17YxSEilF6ApHOtrVoUAjOnf
agqhUTVS5RnLjm2X4FEIKi51GlF+nnk09Hzb2PlABFLh7qP3+P1XtYWCCYxybl1aVSZUtSVQAeXU
ZJhJqovVksmTqn5zKpKUhg9hp7/d5LqefLtUMNa7H/ZrieADsDrt2ERf8eILRJTXlTbZUBD0Ly1n
qAw6KP9SE/T7CR+MyWg+rVGVDxJ6Nup5E1vXOTJtTsqvVUsoOv8uJnIMTC5LRJjM0vqtE8rvxE/l
YIIngcFRGU6/byqqcnoLxgdRdmP83GFK7LEnkLTyr/V7wCwM0MSbEuDsZdCUS/ZuwYyVfc1Sax4S
bRFS4crWaQoEaKAb0SjGoHolthgBTUEKFUGoRMHmLyStmRelIFkmuCh/OuM6XgoMpEdIgeA3hu4O
PP/Zn3W7PN/6OxQ15MZNSkW08hdPcPeefIqiRhwJfIztZeGd76cUd7Be2k4oqCX8yv5tQjXAkqNN
MeRGTLvQ35YD7Xo6pnot8urdrmNMy84fKH9ePHsgkNjzB/Gb5rrp5nhn3f1io6FoAXqAjco93vxu
EEuqkSJigSzrIvMRhkq3QwIbDNEQHOT7EaFLeEnWNWR9m1p7wlDHRRIwqJXh8gikTDT9zao4uykC
OcvOOexn8QZEOsT9AfLsKh1Q8JDVGm1lbTldszavGTwzjdz+yxvbUGJbBcl9Zcg6kmfA5+wkKrle
xJDSRYAP/r09YcWbImaV//Z3l9lOxNCZ1UiCW+awXN7gbgctl3hZlrTgxrHO47Llz9L3QQUPMRVe
prQerl1TEs1LmBjov9YwHvMIK5wnnkVgE/tBKGdn6dn2idLl1MsUznnxOKaOXs1cNwqQr+9EhN20
aNGxiWRkzbg9ccJaLxfJpdUMefCXfj7m2B7c7CBCQWp7RcyKFHSWAxie0c7p1ySUo/787EjV7K8W
n+9xEjMhBHTJ5GQEG90C1fiR8uAiedfTbNiGokD9yvqNOQRBt11fAfisiFSherQRmsCDV6el+7co
28yxVDuxDSYvb8ASXO6pedN4XVmFpnQWKshr3l5NPxS8PZY3nESTXnDsG8mSBZZacU7ucKaXljvh
M8P228j2nsL0FTeJepsTQRclcA6v9pzYATrrpix1rmZ5/uVAgnAkbMe5wQ1BhyLFgCjSzbCdFVeD
0uIANsDA8xoFCKH7EGG/TQKK37Kc1hTsDe1N+YjL4J1h5NeFT2WoWlmgxhUsW7QToMvMzR30p26j
fLnaBsI6CQ/omJWy4qrF5VVhl97r0co+LbuGX4FugG2YOpkYtUxIDadZfk/O+BErtnvFQp7dgAHj
KxZWy1FSl09XVWWL29O30+NogmORYlrSjd4ZEnJymjPWSMGb7Aw2OmshCHBaJkdW7bvoyZ3B+FMw
4fCMgnUOp1w4coIQIsqwIVaWBpl2acJNV9JyN3J+Rvs5CUuYRxBJDf1X1g/kTCZ49UQhdQd3SQjJ
Jag1Z5tX3rkAbgBL+uoEWV5ADMqEiGx8EkoyVGKQaoDXhEqhkd3wlrerraIQ6WK/1VLBlp3Qq2Sp
AB6FRGzEZV79NvYEYNJe+kCS2R4kAUAUYI/zHfBd5KOYBE+oInJWMYTa9R9Aqs0idSUaXxVv6n6w
MRwxf/F1g8c19NIB3UvLF7GTRvOlYI65iYlA3wLmCsQTNJoxUvHDjxyCLmMLnSFbPIqHYzAelq4v
HIF0n/ms7tnG3XXfqD6Jga4hvTiD8mAqgLQLGe1JyV2KcblZlJLgNFu12UwW6fuyAx25fqrIRBYp
/caFUY4DpxOHsWBih3/T50Ktpj658HK+BVW6+lvf22XOKa82cj76EQ3l+DrsvAale46Mosn0vGVX
fgqZ6paAtCsM9wt9ipxlGJu4wkqK6b8rIfMBfwgG4VWO5zxuHgvvrAEDG7V3vmf2jQtETyl9VWbz
ReLR2s+NiDDqgZSpcg3HX5b+Ep3wHZ8VTm/s8tOdms8V4wGarEXzOWb0LigGH382h87tktQZIqNk
2eaMFIVJFV6erJyNfZQJcZpPz5csiRKDg1eQmTZgfeJxwycUM3SSd17Dc/f7mD+vZHrqkKIIPW9O
BIf9kZyyqpibtAd5n2fxDSCZ0YSawqQWP5Gs6mFfIKR6SdzOUTc0/+BwVM9FqcU4AQiP47GrCUU/
1yJrBMEW+eH11tJ1HeMEGFqM2rGhXYVzWOBf6mXcfKszv0mUxt3igbAC+exgWEP37vag3ABhhWTu
/52vJx4INIAN7rAF51vshrqwc83ggI2e97nS7AuECet0KO+0EJnFwdLGDI3V0oU9ABqGoP8Q5LmI
mreaDj600FmJojcBV+TRol7zqKHKWcaewH14oiURBXz5rMWxLGHf5IAjIDc/s5HOHjilrcNrdXsJ
mRKS6siXJC1r6eq0lUjKTXEiod7JjYgpusTaXicEFjWx4O6ds1Q1CZjDH4Lzg9Ab66/j2qUWE5Sd
LHY2rxmgTRASh1fmApX2WvVDWT83RZ6A5lPCVV3T4N9hNXmgEfSU54c41bcn4j3VQvV4729oKwEM
4ZL2o9uTFg6j4MWinpRpJqX5xWQ5bP/sUwzAjYaVIaGqr0RZUuxKTVuH8cmI7aDSTMA0SEqH3i++
7by9XLMbewqG2oEZLZA2LCd5azqkqBhsyDlKoRbOeIfHBA/FGQBt4HcwcrqK7HCyRtdh+JaNI7KG
xyu5/1vGQmy4L6zRStS4FfsUicwegAtZNWveTY6u8XPeFLzC2pw/UXHSQgs7YyKImaIEvlmyHfCp
9NxiMGWUJooq1Mkaf5ShGWZD1EGOMzt9OVnkbBW9n5/Uq4LeCT8HyrS3kaGPJp5IsPWrAg1ucuRM
3wwysfFvwniFbns+6i6lEGV4QZg+a3fIGVNskSEumSIogfZjrks8PCnAGy36pyzqgZj//Kws5CdB
LlXDdh6fwFf6lOVlcMlhVBCawoweUbyeLc7XbD+7YTHmLl1l5xAgUiJeEvXjDEeeu785vUt4KoX7
OThnTCU1z8yX+0hAZUd+QdFuOMG8AHDadLRffc/tbMzaE4L0npDGkVWpY3FHTU2cYwn86U7ScuDH
i2LcNUBOxNdMB9wFODmutTC6PY0v3vUO8QlFHPvyK9nkD4ZbmWqARRvti/VYa4KXrYPigrLEA+YP
k6TvFIayNOrYiHc5cxj6U8GmWPibtq9jUiqaTgUNeB/h+dUBRs5pI5+a7sfWF0IyMNa/03kKrk6v
+3AVesRYJXFQxN9Cth8bpuOI9F9h0jr5YBBR1ipH3OtCUWC+SOcji/+reKtyu/DDToQ6HW/JM4T9
KuDUz7UugFV38QnMoRh9C40ivuAvF0VGcXh7bebl9Slid4LK+YwGS+j4KqdNg1hJrKHCMFWG1sX0
/5Y8v6Lehrqu0UAJC/A2e+eHM1+jM16VrsperXcvV/uejy/4dljrKPUO5rRJgDUHvy87Qjc1xR3L
CoxQ4hQR50ZY7K8C+ZszGcSbXwTkBQfGYv1fHd7hRjK8ltnWwRbGE4c13vWL0VSxtTBtwmu2DIHp
4f/h0MuzR4hD7s7mcAz0tYdX0SM7zjjH7DKCmHnnjnYLIl/BtwRE1P9OfaGW0vSF+b/5YDERaXYp
vbZjk0PhkRJszp3skAmzr0XvA3GONOeMELZWDFyZNcD3IXHWIP6bJJ9mvfitDN0GvmyhFnSRix57
ueRmORkRgi9Z2A1rRvPzxeL9zBD85wGHrZQbpAXw1ZoBntVgpnt2vTGF9YLjmvwdvC+TJar0FkIf
WHtjTw/mLnQ7LR5vF/NXcW79sAd/zeeBST5x2eQtZhY5n2ujSvybDn1/vhfNOA8LnQjmJzUUBqzg
EtvT1Zn57bIMYhoa4D3gGbDe4vyod5qYixgqzs5aD8v/cobCohVJnb15djyYwmCgdmY0/zbQ53Bj
7Bef3bBZFvcQYFGnzHB+XZhXscYICwik/1R8+IBGPi8sZjQstkXcN2Pwtch/+8NbuD/DT6yEjIFL
QDbtSilRXCyMQH89hisbzAtacNt73WtEJ/igWT1AXLiJduB+2z3hwhWKXwtkSiwn0gmIcAxO8eeP
iYOcsfqBcPAn8vfbAJPVYD9M3sYIi6YEGaIHMUhaVB8RswNk79xV2DYmt0XlCpiAo1YexzMZaJIZ
So3ZcUScDecvkaCjEH7p+VxNm04grM18KLNVBRoFDnn2E5T4+ahhjmOcHBGC/ffsRAjchLlfyHQu
Uz/2N967XpAfVBEqft2wxBAc3LxNv879euKGpU9gxYgBAAnqPZpmMFMtytTALwc/dEFtLw+8Iayp
z+t0BQ4OQ/KxKT74xSLkS6Ms316oewHBNTiu4fdEFW4CUN0oWC5Gj4sbWRhzCbvWL5HtagD1iYVc
jUXCXLHGxOZxi9Sz8rHUhodxCgw7Zm2bB5D5BoVPPJ62+do+may/EHwlshpVTJHRqRgWb7y9J6TQ
GXCoUOVIRXSZTMM2mT5dKOXXrFmtO0Z110wLSlwlEygUDAWC660DRs2ZQnrF+O28WcOZEXXBL/Jh
tHgxeJJnfZGwV3KrO48594dqvFrJOQtv7SDAF7uPlTa77QJTrP2Df/nhpNd8YpaudfcfeukICmYw
dJhFgU/XbbgnSzlN//L2UqGfHhQurDV5XUsI9+2Cfk684HKFvPhohEoK5FgrqAX3PP3IumOGxZWJ
hP4Azmas8KIfkYSv5pzneiOLRtAyRONaH4oGobbjZoPIBB4vd01gHXqu0yfYChbe5G1uUVyyWyGG
PmIWm89uo7w/gtpXbF1zb5lujF+jZt4Qasbhol7El2JwsaUoNEwlYTnuYLV9+gwjCjLOvTEYwt4x
qK95MB6wL/ChS52vChp9ChfFiMBtGINydnKk9nCGkryvUiF1O/UqHIJgTXhhCm/NwvqZ2KniXWiH
5BVVgG5T0WcWYp1x/cyNEOuYYfZ9kk524EU0BuN1EJb+mFWQZVTX+f6/DzaQODD0F582F7Edkcar
/aT88PK9An5Zrll+e4/mPXGFymwgITJl8SNAa21GhcS5ncZzZ8ckw7pZiZAxBOQHn8DObsyqMRzf
br+zBiDY1TBjPcFF1pY5Cdl/jpSVixkLUeTDNPiIR/M8PkY4KnFZnlYc8miCm6u7aC4MWK2F9wH6
nIPyEqmdyZfVos+80dBL+Z5PpGuIAd1TU0Y8gqWD8qtO++kcK9v228E/KxIkuDKkMCF6IGn1QejO
9kJ8zZbdvgJQz5qTsbf8zdXWFlV3jOQ8jcGAPUCMdTC+HkBnYf2FTsYytFK/d7wipxSKOHt3dMTF
ImRa8hxZoj4m6+2mZ1mjgH7XijuD253sFh3rwJyah3EdbFn4mTNb5Dy1j30W1ieCQIhhJDaBe9PM
nTfK0US0BMGTv3uYBpScVaQElVjkJq35Pd7bDgAglaRgDwzxO8yKAO9cCHW+3NT88fWEYAJJdhiJ
9gErT3Si+p6nPudHQDomRMTDDJa4I3UhZi5FJGihmWXPRoUrDlbISWlbIrPorr11GXHz8Xcsump7
SMEnM9/cyu5ccLC3jw+On3ASnCsLHnB/Ia9esPgRv6NiQl6oDsPt7ng5ZpIYOsUeCecSAVzNmugb
Qsz2o7eups0/ochuv/yvS9OGZcnDiOiatzXxOkbSX6Ofkalyrn/RhVmYH7HdjyMOf5ROpFfpcC3Q
8CcdEOQtoj8lxU/XyCF/aWxiG+RPsOa+CRe/Ip7fcyrbRBoWn0fcEvKNFYscRW0O8YVNggfcT1qW
prMAjA8w3HqA4uIe2NtraxiKSPJjILieW9oc671ZFJ9y7lTLgp0/lla89Osk01bf5sIB078PCi36
umKaHJB//wfNvGHazzXm3I8ORBSsmJa+s8TE7uoBPqQ52Y8/sGctA0ApQ81wpBiZwJkScAELs2Bg
+bVNoW3hOU6ZvYCCaILa9vYyUBxPSRDczjcV1HERD1fwgaG+ds9bO02+35dkBCl3S+6tIRKxGrRq
mbfft0gOMLx3sBsfpQkV1bO4pz3OA/wJfdrNsT/G6ByfwmunX+G+B/xjgASHf8goUNB0+EmijW5k
eBr44hXt/NZcvEOj9pba68GDynP0C3mC8hhOI7Nrz+HSVxPJHp14gD4NFRrRV5E7M1Q/YWqspdR6
jGX7JC94ERb6e/84eOeGuDBpPqjvoaOMvPPC9lyZYUYnB/T8CXfHPEYges+2racpr2+MIGIaqRm7
QGL75Rw60vUNW2wrRCLPCmimYYgnvjajSp7lY7Fehb2EPTFU+WLlutPDAhay9rM89W9w85/hYoHF
LoNfyR0/QeoEQAPcTLMyb7sPGq8vn3pStALH2NxHNtZ38EK+OaqZfs+bgQ32IENgtLcXAf2rf0Km
Hbx/3+vInEw+Uz4KRNO4/HSAMhA3fB/NpNJ0/gCL8aJ2aGlIn9HuBYJRMVrgT1v92HXNQXdpfv9Y
KbmAjZDIiubR6jxFUj7dYl+ZNrV63DNfJUKLYn6f3dwnoNKmbzSYbhTkN8T/+EvcZ1kQvrH4WkJS
OYkd/YMeLZAMSNK5WFCpCTBMtbXwcIPS8QywAC8NKMbgDC8dcIUpCV+dwnCuc3jQKCYDJkd6iPZA
1heM2ADt+ZlnXh0U6RosGXh92qE6bKMGs9U/18IKd8l9gfq7FahXK4qCZ55SNSTejLmPCT41IjC2
1wycMaL3cxePf8zWyxi/SoyRfKZDhOsr8RZt5kTMZ3zBq00scQe6TltwSI7OlGVHEracFJGYWSYJ
KJiuRxNQr+EpYWRp0dIf+kJIluGNhUEdTF2AibzOam1xZwi6i7ntOGJIErcNbxx7y6nUiaLItfXc
69AEzIb5lWUd+Rsx2MCrmob+JV0NdtL7Hr+zYB0TR3ldBEJGJxg4tULW0Zyh8mMLXc5hhEiN26+a
pMk12nY3/7eik100cmoWa04R+Q3Cx8FfCsPIh7duCnElFb5cZT1oXvCy7z6DHqzFDh4ZunuozZFc
wVXvYwtnw9Lc9Di9e6ysd4jJZN5v6jSXD/navIpafc7VF9CoJ5+bYYL6NNdmeNPhiq+29+iEhGqT
73/H34Zu7ayJDRt++2/lmN6pLwpOjR32vVg8IwXdUQrSqQju9VdFoMEokViA8VUCQvKmkeTFDufU
4LW736Y87pmZhGK7Gckq6yFFN3TW0SlaVB3da6VV3ogGZCiXznuw7RiFWFnFTVIj3V6fBmOY337V
oPug471yi3SqokQT71BOnvTOHPbKkB2bxnHKmF96pdBpC2SAJ7wy9aRNbgvlzDAvOlv8UjsTpjV4
/PgDTHPgt7ayg0WDX2wwwkmsgi7Um+ovl6/MO9qbT3m8Kb7zXHTMl6jRDz9PV58tSirQI4EcmtOs
9m3wJj5y+/s6ZIvanUL1/rodxf95T+W5p3SIUsSoHX1U11Sv3/4KSCgdhITMEIXVkb/y+WNxo88b
noO5BK8gEF8iSwjiiVRh06l9wiEFpfxmcQrYvSHfZ3PEyHgGjKdD2xWCxzcIw2RL3pZsJEKiB5hg
d2b3L7m0sfqa5RHh7U2fHD5kZaHJYJL3a3OOEMXgJJffDmrAV1QSl7d8K6to3UcnWhTIEOAtywW3
GouupJac31F7e+TXiNnyZLQ0OFF1XSawzrGUSal2PmPtHuYnRbG42zBXJsOTfCwSqvUFpqZBD4UP
Se9/gD31c1AKlcKBW+Pqsa0NmKAO/HNjQ8xLgqSauvPJE4EW92z5GRyZJpw/Sz0SBlt/D8WYCN4j
njTVQi4x/5CQ6w5tGwUf90W36eH1OPkJF9SpQf/hUnFZxYsAcNCR2rd+TOfp7nFktF/PgEI/O49H
seAt8TIOfJ0rUX7rUVQeR08FPydvoRDOwX+HrPFd34Yr+W+O8cJYYDBVv4pja4WK6y33Ojhj4dYi
SnaJGFnQtYbxXpHjvCo+0sv+i17zRwvrW0euCROci7vexGktRrWsoxuB0lhr7FWwIgM33xNxNBoC
cJoy25ASCgelinSaI/bHi5lbYdetWd75BS2rAXTP/QLc79WYTvWvGDO2JIXFFDVaSpp7gOnBzDtT
U6ytt51ZUYNY/df2C+N7khbjLJYCKY2DAeRjartm0KQJjrYu93WKr9hTvV6oBEDYYVtzhz8s4+mR
5oNrgtIKXzZ5HI8VYkH9vjdXnji2dpXRXS/vFiItUkK5eZs2qIsBJSAwdrjkjdQy5U+CGp5FDG4Y
baOx2BzB7UMQUyNSExsjImrKyoFnG/VvfCtOo6eb01UoWoImAkQgu3rUI4GpbkTtJ0dxj6lR+Bwl
IXFumtQmn7gIBtYaRuDOeOvDdsTpElu5b1/gHT1fmPVJ6DnzXWq2gpkKITsuM2TKfDRZ6zE6td08
vy2KoOJ750E97T5if4S9bR0br2icQIt5xKI25B6fVqXYvcd+Ll1k12089XeJzCKy3eZZZGlNxNk2
A+vYDabd2SfC1f3cFXAt0C4s0qaCrDXB2YpuM1YSf8WwhSyatrGUAX/ePK72djqhwOfDCjjE7gNH
YG7GcwDQ073fP9OhE6BpAO9/8YtsLQgG2mhcp5HwktvUa7QZGuJigCnQM3ixP9AkjWvsJtK67/KQ
zQx5JqWbeQEc5+cAF1l14qGfFx/0qPo5r+a5r4UEwEXZJ/kKYM+wtqqUncB8vPWTbYL62z69sHVE
GaRiotsUqbt8W5FdgiHVYh0MCMZ/086V++uruOIBNXPl6/h6RfNBmuJl+TFOa9OAK58NqLObayjn
nCV0r0/GM3hixVCaMv69n3PR6NCGYOOVHZ7Tm1AFVQBEeLliiAqS0Pc9Xu8AAE5kfDQ6aWBBwu0P
ZZ7MLH5OGMlDhurD/EjKbqtl/77QQ+JmL48ocMdSu+zlVm/2+f6YDdG4rXOjAamjNS8PGie0IDE0
YwspOPudYwaN9cYLCrhcdsSoCjFGBIJUWBr334yV620TAkTZFhjMVJVL4jFnOH3CvXGJDCFMjLbz
w/T96LFHGjLuQ2JFsU7RMcVsKU/z44c8kDxgj6yfJ0CyR0S2B3K5LaiX9DEJjqYpGhj+PPLQ/J8o
c4Mg3Ndo/p8QBl1DIhO2F+1NZQhFy/YdC6m7K1Vo7goo+sC0xyCJ7XZVDa5tOSJA91KsvVB0X5e4
kQwWumTpa8cF2GVocPyQojCWwNtc/Q2Z28a/x2a+5C8CZKTR4jPQIIAod7fSSP06Tlq0L6yPd0lz
gkjtehQQZkuFu62GHPjR3Em4PZFN51Tq1jLW6BlUelAJJ1YZm7Cu8/F4Xv2i8HKNQg8MTU6Byzh/
Ix9tah9oiOlJKsVbVwcD5Crny8b0zLfJnMO8SZo0ahkDa2Ie/saY4ecG4Cm/RTT5HWuRQicJWp6e
1cF333EwTY24GNrL7kOh5CQ3sjz/d1fL9C7zPSpIZp6NlQd+WtQ9aFlFf+y3PJb+vVkUf1thM1fd
Rtpc2//zwhnlJ0bEW3Q/kcGydptOGwOWAsFq9bSdNcAr7MhJ1HseO8cQXEK77r14cBgcNWe/Qy2K
utbKhYA9657F/pxZpe2+Fnx+YrYvnAZcjLzJdnzK5blz8loyxSMj6j2H/xW/EbKrr3VH81LF6PwI
sYsyKhbiuWu4pZ64773FJF4anLVeU6OOlr1Kn46wpPyh4q6aDkgq/YZISV2A2bzxr002pCcwwP7q
rYmuNNN2xt0eXQEvd64VjLoOXSghHdOAxRAAxXnWKvMkoV4xOfdJAGFaempL/sP+0+tf9JozwasK
5dhdODSVTqZfZJQoprJr2Vk+6T5cwvHiLEARMY0zKjrL0MNp+ET1OF83QUjay4YoNK6TXZpvIBEl
9YfIfqMTvRJEOj8/Xu9py8MKgOUqpabiSgpWdKoo1fxaTqhhDCIGVmtQJug7BAYsc2rnnM7rg5Nb
10UpM+MVHzDsicQ50TBJillL6u+R62NfynaXXJDGfojDL2B22uhRRHQsdQLOkTuqvxHyVG3MbRnu
LadYDF2Q50SuL6AcveO5KAq4sbf1nOFjfi2zlmB8XobNN786nvRQTILC7wPMKUJ/wEIow+u/Rfiv
oPJp8ysFzYLUz2ZBfB8rjZvIJYKz79cxji+lRVE6gFq+IKVcOfjqd5ABDEj12p0tU1Dond+J8iOG
JYJEo1JmSejJz1WrbtOY8VJbzY7Wef9r/5biebfAbR78V+CSNMI/Ps5J+tZBN7jbl69ycQ/NXeFp
QXSmMoIn4Odu2Rh+Pf/d48MuzoLZQkpG6u/Rk25pQGIZY1ck+Qwr0w54W6Nh4eIyromjp5Ko9k7P
e4f682WHCpb3vXB8WQAt/fRk7Wq75Mo5kPrkzdMA/5+E9WxIRQBAPtNf8Wc5O5pLXwWh4G0BB/SC
Tx6Ufcf3qgEhfz92vMr+DklY5pakLtDeGRlSfqWYddNncHCeeGV//wYxmzT9JGnkOR/pjmryC45M
1vLeq4aws49bM6DG+XfFjxypMPUWxwVh9ZKzXHEfdZ4lKFBV5fe09vePzXEjWZRDd/VMd+R7ohbJ
DJdmX3GJ0CZowIEKvSkfsEwSMFomzlT5VDzpBNiMQRB7aV1Jjk+7f+Ft8PPlvM40lY3Xtu69Xq6s
oH4s/pJFO0xEuhtXZtoNUrz5TojvgsYJzTAs0b1vYlzxe2GSVXo/rEY8tqgPbrTMyP1C9B9BlpXR
swfwSyvcckgEgF1UIXl7qoYNMSFD4UFIpXrkWoqI87/1ZWEfJPw6rt1DjKEl0R/YKkDkkNwkGI0N
ZtM34uDK3UrNldRlRQW6+HBvRnPtwAVF+gUhER2E8o1hnd1wfyhCYCE4WSFCBVVmBG/6H2ftADUn
Fe6MNA2A1O2JRZX92Q54XVjOxUbAZk180O7sexKpx1CWoC+zLpoV+/9Ollnj1eK/K9+hPu7zJJUO
dRpO5Y1BZV55Z7m2ezrzHpN8wrv5KATfmkhxnDNRJiTf9Z0xuemCrjTJUr11z67IQdw/NGUXiHm2
FfNrCr4ICmFhts12rPp3Qb9lHrndGr8xD9E3cKmrBSlNF0jcMhX0N59X6csQZ0Y3nCrWoS4PazMK
tTL8mhxcnx6Op0XllYogfmBTmQdugQzoXW1qBirA3IZ8/uSztOKDo5Os9u+h6tiBo18Q4jrKzmsC
OmWPQ0I47Bck5Z6Eajf8M+muDUTkLTM7uA3IaaxMgnAEtX5WMa23aAbs1t+Jy+oB7i3yDNFGduBr
k783Pm/ViYu2YwgMgTxnZHstOz+qe4/WAW780pwhh5KohJFyoMhGFhyP7cCEN80gftPJfIMhDjHw
MBWQVtnL8Y6oc344U8cnfIYBMt9k4JcOfMVU8fFXrtwexiHAJOV1utxXsPTKkKN/ystgpfcenRSC
tynzl46BnmA7Iy4Un3Bqjgl05tABL0SKxnatUTEOOKE0s2QV6WcDTBGccw2KrZqPx/7Ore7wz+El
mMC7JwBv3tPedLGLg148jDvWNiP5OLGbCcMTfc19U/fxkcmvG/f8Ts0TkC21QKIiOg5nN0cx/kHE
KqJJr4hy9GaxXX7lDDGCIiP4cYijJChKfU63iVTS6sLyRT0NkR+2QmagjzU8nttsGCklhZgPBTsr
fnQT39ATIMfo8w0jzmILXcVswILW1E5RQfBaQdl/rh5SgFZrZ/JB5pFSRuy2MX4CuR0+1PLExHCn
UM/XdVLqEHgv7GsrOg/Zl+ovRw2mWJ3p1D63tEUWwt/CreSesdrU3qYbCkzsOEpyncrcgmwFqpd/
MnpKojYAofwKT64C9kMCV3o45u5680SSVdE/aRs7y91K9ysfKpl3646WSiO0R4TEJbqahT8dJWte
W+XG//d8NHu1/ihyMGS5WHpc7k+4G5bg454WvZTWC0p6nZhm8at0sUJ1t74JU0vxKL8nKsbYkhpc
6MXcWwBoCXV5HeMDBGIaGCPOvRs8aB17Doqa3yv28ZDkP/x8ocpYOJW4qCvnN5Nu2iHC82R74nEn
WKcbK9C6+d0vmr6Y9X5y0e9kMUYiaHwioolBCw1g2b9cuZW0+yxl6EwcZYqiDdBbIPJu9qISBAYe
RLlnk2GnS4P4zvxB+nEfubiTLXsv9urkrk03GIADjkayrM4fFnNjiOcpLItlvWkAYu0b0/DpQDte
UrlF+A8HI0OYbSyuQCzWcuzzaII2mJJuFkIdpNz7QfsnKJWvNZVqJF5q7c4QFP/U6oa5r3w+Sx4t
GH+jBGSWsQahgk87yaD/nqxRRY4Rn+cg2fNaVYTRXTN4BeH4Yc/r/9TBfmgrwAZTNR0txV2ACmzr
VKJ2V/XhC4RrF41IeRD1CM6ObC74zyh0p58VKxUXwl70qX4HVu0AzPHEGYrMlJn/rQnrHRzWn9tn
/KYvt4T7otGC8wdYNkm3BY1CRf/YT38jtiEqZx58w7zY6sOiZZ3cshwPkAoHfimYH+Gx5vNkZouH
3g9yyV7atgzH5OQueTNjO3ocNbepswFNr/3N6xZAm9gGXiuAtny8bqWXElETT3n5DnHqjcGPUI3b
8jsnrcj2zQmIA/vzNuzxLmXlA2ljNivj5Vz8w7MI/DLeDHh2NmDpYCplfYoP2cx51EY/+ZmRvHNh
sEEIQ+1ZOzq3PfgxbbL58mcTai6w2vTVZuCnr1ezCeVDa8w9zWvsox2do0fWoUK6y/h6u7EICyWJ
ND33M82/9dOJEbSUL80ZF+qhOXBCMT//u88Fbulc9tV9FtD9Fc+0jvjiCgp0nqSuoFk9zs4nVdGR
n7l2tTmF2PETYJ5Qd/obmdHSGSpYtUJrcpZZ4GuOtlYsizJNs01LWqgH1ebWYpMOeCxtzm03EYqb
W7o3hZSLrUiNBJ8qRvk2PXLPsfNsQnc6LSiLkLsaP5v60ouayES1K3jlsQolwvNcqR2IV6/VfnIV
rCWvPJr0ajpWGIDQvry0our8HQpnGR7Ts65fI9uFIZP6ZYoqPRfUG6idar7YTAu8vaezYPOdMlyB
cVp1JPGJ+Y+Vid/TzbPurHM5fFIB+euLB5vjWmpTsQZ71sf6n3fvs49dPKT0Xlc9cTb7D+CtP6vD
o2eesClGRwFpIur8uVc2feW76UByYjkR51YoFZeZ4G47CqyQ1kFkIPxkgnF+xAAHe3L7Un8SfrAw
Q7zUyqDP0T1egXKn8vitdi+OmqqvYMeJvAmv04jDpa3lCEq5WagBuc3BAhcc5QVpP4hNXmkJT0el
1P6xkfwJJh8FbzcaYllp7pVp4oEVTePQWB+XaEVJ6EP4/8ThKvfcEjlzfLlFBnOTJs4gnqmoRXWI
wulc0umjUbsB5lgryGgAttKEmR4pveojIMa3V5ExdkFA0ztCAJqJ04gaqGuUULi0Psi2KBTxZM04
ujCgFTXpyLe3HdiM5geHyPTK/kWifIcBb7P7S1iKX55vZz0CKgHJRcMEOkww8hZ2oFzK7GmAdfID
AKPA202Qgm5Z175m/SIVGGfGitSXHeMDddQvsknh/EfS/VW3Nr+dm0GuJkgKgLWjzLH/TVHfD9v6
vQFKvA6td+BbGvig3Q0mQKgV6t9D1pe3S63zxYox0K3u65o2wSohhI4OBit9JeGKB99bWHctDtZO
EJYFbREI733Fdi2nzw4jrAxcUbO7l2yF0torBfaNC5j1eeixtqtHm0fq/IGqPVKuaRp+9ImjG0AC
VjlB93tPIfdxiEe7n60EBmqneSqCYt7+svi6HC0tMwBFqAeywgUKN1mBjgxa4Ju42cCdhBk5s3Xz
jgWXQ8KUzxGPlDrAMR9c5Zdbub67uFR1evtxew4hTDYLGEwh+8mmnyzYGMbJUxyo0pVWehhZSdgP
jmqQjeLskk+sbEwdxYYR2iPRq58wZEm2FTGrZdzjGaE9AkY+Cx1f52fS+uDnOjnSALZFZOFi3e4+
3Qqg/OocXYmhx4fM5xQ02HlwEO3oUoHI5RKfyP28zGCDyrp6vxfsNlO/nG2YUwwGXCg+iY01uZIx
bxijE3De2YhETK7DjK3OA8k/OfmU0SoS1jR531colHObUZKcA1L9Bguphwh0Xc6XlpzBZVtTEFj5
71+Qe8cQL48py/xz0wieTWjLXcoKR63Rpkl2H5yJUoCmcY/pdCgJwH2CD2QTHWGOvbObKHS9W/Ab
hA0VqvKtajawTRHL5BZm34UZLlcOInQE9q2u8DmBHVxPqNvs4RV87C0VnSs6k8YyPLxq4x26HCwC
rwsgnlevqekPuuRpVOj+Ay8AXMUxnsBbV1pZZtfdbMHBuX4fMbttup9/Kds3120k+qPsK5+Tj4SO
ITFsjBZaSEryO2mizTGFAXHDHy/6irLinJenrKFfAgPU//GEbJBgqGViCCT5Y6ittVbgKMFGixHT
qt569G7HMcFn0UdemEYlz7+Nhx1jAhDsGd9OyUBrfL/CxWVnhl+fU43tx0n6Sdbt3OtF99HGz2qe
j4LXaBpCTFDdaqmzDWXqdMdCEKfT8WljnbMsFV746hyBe9N+bINH4gudq3G4Tx9P9hZs7W5n5zgd
fHluGMFW9VPC4XbyH/8YmXWwfBYbBlccwS2+LCe16NBsis0NNm++90hLxoO3rn56qyiKQ0M16dqs
jkp//u4sLNdo5j7CzqUfpxMikoGwLgIu7OuphM22pALCbLK99QjSqjy1mN+4vl6cC6TUZzFe+ohQ
0Db+MCT6nmXIW/Ll4jXNBnWV3w1fRWWeSE7OYVQyGqvWPlQ8+RtQUnhHtUfJjgA6oh+Sp6sam6/8
RqkRif7QyRQQKpcuMsxA5k3Ug43bfygg3zyUkDFftBuJloY8csC/tqQYQbMw3apUscg12amr9Z5+
MDrFTBdfvd2nPav+g/DnMTGLOVa5TGN+NhIdyj82YKnrmBLq2HjvFfhsJ/ejEF+w/7hZnAFodz7q
XZqM+Ci9GKI/FZAj0xV5L7GfcTg3uBqR7aPhkiz0N0vXnMtam2fdZi1QkMUteTFzyvVEQAGI07qj
OcINne+kYDiQwyOAjNlpeRpF1Tm/30n3mhGtcCEyMIHY/+5GYuS3/KF8Nvaxv5PumjVeiaU+lU9t
r90P5QSdCBzJMpbpECjwTGNoIB/j+gasF3VdEjfkghYxmLiD7zA4olBdMXAVtL8gB++SFJTAXurf
cM5NC4hu39wOz+HEMpa1l56c14MDzRKg4//xCTGzwy6kA7nLnHb3JpxiPvUu2t41w9QmWzi7oq8E
oGIrMdbMYbE7x4Ei1RX96KneO+j+uyTSlI05DIT9X8BfUnoefn5G0wMM9w/HFFnofVsQVYU3uSJ/
8PTBsm0rPC/3bjZcisUAZrT9qAW8WsA7Z56XDOhciQJZiEqi9vp1LwquxdwVaqVVN+ncpkg39I9N
6rBXgX/ohat3SoFhOR2RHW+nL08SMvQU14c0gzGu3T5kzKZdUdvn+NE0RKrr1lkO+NJwYu16Yr8q
Gc2DvzRduF1ic5COm6cNaR0X0rEN1iW7mqNg/rgWntgDHdj7Lhk/mFle1+WJxcs53smwlxLYqyoD
xEimkF/zD/cGIQnB31M3pPILQQIGnGwKbXyguzVueu7dVXdniA22Sf3fXIaPz6FYGxjTY0Yta40Z
fYna7QAB7SQCs/D52wBplgDu0gUwCVaMwD33t2dpDG+QgJe3nNTs4tKTk/zmyq0vD1KevzhHn+N3
l0yWIZpVzhoqa6XiryihSv2a/frKGOdsZ1JfCYOwBqQ/D6ZqES6ehDqdMflxkvFJBC2LVM4/o3TH
Dol66v7i0jynoHjBodm58stVXfXAUL0TRnF3k0peKyy+ZTaOWDWLIgBqZTRtfTh//bjdNhaDs5tB
9O6jkrz4wGAEH2tHpb8M/OY+2DjCJ9FecP5zMmLYhn7nph7I8ThYWG3hTe3LHTie3QDeydo7s8xw
uBGGvQonc6NX5Y5z9MyV9/sn2Th2RcoxJDsw0Cmv4HE4cFoyi8X1GpkWiR5iyAgFP2ASmfrDq2fw
/vRa0q0Qvmc/EEdgmxFMtfpHVGAtnYklkoAZZDQZkQ1PiLvGuX/57+MOYPCgc6rWYqOGhtfAFQHD
fjxMe73lxCoTxVti7yCGeT+dBDXVjaJqNUh1twfehWPInaPg6NQiCPerN6JbDZR9M9ji9Zj+6c5D
mMMOD3lj5GBkxDOOLAuvmD635gLm4gm6N+g6i47yR1oA875dRBJ5jKDCBQNEF4YuZTlUCp4erq8Y
TQ98gcCcfYxDSfiTOwnJs0WOAqYfAT3zQxOpZD7M3Crmn6/ljOE3vBbasRsgAXzvzbR+rA7RzS/b
2kiMb8w5vKymKZhtgrThIFY7baNlclktsCO2c6IJoR5CJmsK4DoAoc4DbVYNfUSkxB2n4b38GO82
EF+gvCuMG+6BXcnf69dBmeDGdc6RsEMPeQZ4GWNHfBStCCxCAGk+dqpGlR+DhA1ercez9bCVaCev
NrgaEWsnHpGjnLQTd53ydf3+QnxNppQ24GYiQcZ7nxH7zRTDlyHlOTP9pGG8asCkbRd0nMNhgK6v
eM9jnxdAlcmpIxvrMynXotzeFl5Lk4RRZgnHH3H9BJcAXA/wE8XsRuLCs4O2DYVvyA8tfs/xWQjz
92J5X0XaRHBOk3ur1ad89ZfViSFGvepu2zW9Lkw65umAFzzrNCxrMyuvBRbBxvEamAMG4/+6KS9i
rXFgxbLoIBRukd+OYc+HbmxpBczk6V8uaamJvem1z3rtdt1LKUhSv6ie6OGjwGT3DsFHTpIolW5q
f4HIldgCvX9LEsDzNJHfqj2OZ9LO80+Ag2xw5UleTrDyPWbMCf/nuZoTFL9ca0wg2DNHTx4okvIF
VRLXegWg7ve31E/tvIR6CAZLxDBRRK19JVTe5WES5tc7AAlQkR1QhAqDRIpfRaQeQHnknCUwJ6gH
ayjCzW4elnT31JzjR5HNWjvOHNzXuxLI0W75NkazTpzydLoCQXdHKIJFSsiiDxJyNq3fFKo7PMgO
76wyWJuVXZxHE9XXjyN0jxL+g9xcSjK0CbG5Sgmkb2LMESNXWGuvAkiSBbszyTYlrINCnLgDFsE/
TYlNZnzKejsZZ3wTY/hiXHmBZnmi0McgZrdS9fJjhM7S9/8rSx01oKIYWQbrwJtHl6zdfEAVuJjB
1unO+zMujr/c6CAlhPyG0JrEZmbfUZEA+H2MqEN1jp7SpxiEJcTR/aBIh/yvuSFQ+j67c4nPbyFe
nzuvWHO8m8MuK7qZDkn8cNuBKhEmjvxLQhpRbF0ZHOdmhOBXrUqmtGyAFLn4jsIBXJLVz1N5mxUp
Z0KhvV3e6Zp659F1ZXNXS7NNcDUcpPlZssfFxMQ0znzZLWtjkEEhEeNs46lR/dVD2FfvTevKUvOS
rmeZDnzLD47O0JdVzaxIRtXtA3qE0JfTDO6Ndx4xo6XCmVocwauicILBphVmwClLwQvS3yKWVU3U
d9U1X0hSaJ8ZrNwILrcuVCAmI/F+KMAns9TZWtNmimk9wMsufDgAJLS9EeaVollHp2SlH20GZtN0
29jwZHDLJ38dgZTcO1cA32vAUueXjE2B7V6MSWAGxtTB2J96JEIKLA+KkuDth/PFn4c9LN1K9xUU
B0mSDjQQYRe5gr97nNIofY33MbujW8uvyd3ZHiXh2TbkbH5v6EOgCiVHWra+/8mYMrzkiOjgQopW
EYMVS62sSZ7UJWCXcMDxUKmntvbDTLx0fiJUQ9rVVwUAVUxIqIEFbeMV6srQAqi/ph4W74MLhRU8
xXVmbdKkAyVugqHHLVpOfbuSXsJTS0e+fxCeL+B9nssMy46AjI3c+IEl6QZnbvn/4JaJZVPD4Xa7
vKwH3TjB0sHMnYc2tP53tD5PpBegYpo2WUX+iKjFCH4IXftXKg1sjRmUVpQCW6JTCt1tnDk+LsrL
aoR9DbUBHA+tc0NFOftWPArftCYeTIObPOGGG6NLMV4Lq/IMCFpqrSFG4wDs/LAfoc+35MHvW742
QRs2fblniHQiqUIW9y8GjycG6N2VyHj6iGXwx/4NYvq1IFLH4VuSOloFYYtGxb9wcLdeUhDffOIA
u1o3uNRrunXaaTq0uSnSvN6czhwTPnvDLBzbsFPc+7CTuuDVNKc4SVG3rRHOFrCJNgYZQinhtxX4
fPSjNYg7AwW36f+jKz7U3sfGY2vdE70AeFjvjpZqXpg90Dw697+Mgbia/QG+hpdaZTWpVUL4Uvhy
t8h74a4lIIme89deBfYCQN25adGm4EPHGwyg7iy+z83NhINJpUKGK/cYaRNtNlg4AEyDp9YE5LAq
EtnuYwLEaokDk0DwJ6bqR033nbNPGV6sC/yXWNYm9zVOyIGm0fZXlGjfqAjlDy+D17bB+7z50FpN
qchdvMIG1WWUravoB7mUnFMmIWkrh7/+5Z2nbF7bdmQIUT/lxOH6W49gX43q10UmVhq3v7oGRHg2
xESLjGlhPz4bJFsg4w0kFP2fjr0z/TsWaxe4L9Pq0mGqQu69a5AzaPDpxlFYO1f3PfufavRPrn6g
g/7qK8IfsuCQPzttYAM1LHeEKe2nnpJIhaBnGoz8ia5QtTOMXlvenakeObZ4224Y5uDVQeA11Utg
pBedI8SELPtH4Ue3lW8O+Jky8G0ymYSV3XlyVB0DwYlgFHXat21PfneCFjEnUBcuzWaJCqh2Boso
4ZGjaUhaQnJKJeqqy2G6fXOgfXMxgBflBGWlL+Zfbn6EbfUeyNh/4sDnbLntYpdPpoSgfe39Pxnb
QTQL3veRgo0OYImtAtB6RswAqUJL6hhPHJJpFXVoCOd0uoeMTxNizau7nklU+mlpd24ITv/GQS2w
ETiJtJ6MuDW11FMxN1T4OS/08+UwBO3Tdz6i5iTy7XeI/OoAysVQ57Dwn0cdVxo2aA33qCUB3Kk4
GtT78UQ+ASTcz8H6QKs/FTuIgqTUerTEPP5BPmO7wcC3hOhEwjKs13zgH7pdxQZJdn1G+236nb3a
yTv8ypssyhU9zKp8p3ppeNRj8yYXN71E0GTXuYeOMachO2hlnXict/P0d0SQUr0/UAtz8nrVxQlQ
biEReMrXW+uiC6ETJo/qd4GEVet6ceYO1U5Dj9gKQB5GfFY7EGHdawUaifFozMIY/XzRhP0VKagi
Yhedjf3sYO/49XhCADzvUHOaOXVQjza/uJFLHf2uTo/nPZ86NKQJbh0gzTwQaxMr18jI6qLT9mYn
QBWl9jkAfKNqAN/dTVUYCc8kseyME7B+bn678fOPhZznTXd0rJMFn9MP4OaygNuXA+5WhcMF2fV2
gjx3PYNMWU7zcJpTHInZO7MvT7GPvu9NMWHZTbwj7lOnWdayFw5KH/0jfBugIWD8tuJZayJgMijB
EQAQFAPmRxvm2TdeGtDydrTUucuoVkbwFPmmJoSJFDVYO9RbTJbIELEuIU63Ff56V++vg4eAkaWG
3oFXHQ5VBsAF8RHNuZ+TcynjWaPw5t4GD+8etPVoJ5NOCS6ytoW7eqPWEqiSJv1w6mXyT07NyOxh
EoRjWqLeSMvdFDQP3N/+zepNUBPhywoXYzRcKYXUkru0+N8zytU0l2oOtb9ILD7TT/71lKm+mUtR
nvYo6AJoNeyYTMYM6ggJlw1yPR05O0DJ6SuYZkH1JC3I+HpzzyOIexFiPQeEDIc91YMDpeagU6M1
mtlM8GvnJ5c6ZvZtDATe6P/X14vQyK1nam6Eobdp2VB+9pmCsg3LB4fGkAP3ehWLacwdgpTKw9O/
72OuLMbUzd1LlVfXmgDwLBVP3IztUwLUmrSTRmE664zS1gjCPb/f17TzwTOgs1j8dBvw77rXudN3
Gx/TvJ7aZGRjce4DlQGR4Y4D8ehr6cND2wx8rrT6WPMwjudKhPnfXbjbPqK4qFoPf6EC9O2mWqij
3FQIS7qV+IT01OHrVu8PO/ZPTistNkaCP9btDIdWKSxp/Vpl9+UX2spI5MsGHhto4d8Cnd78V2+8
vejmEMqbcTh+pAlWBNLEeLu0w2Ug9Kv1yRS83VWun2dhcesGxeSaiZUPTcSE/OGimvbpDhKgXRhB
KJ3WLxPmr2DSsTuz0oPciwbqzlH1VKu9fLJ5Mi1loLvncNJJ83DDQoMB9W65xm1zdKCzlOEeM6Lx
rf3eQQO8A85s6VJ75w7jucxBxDSp1jnrfHwJ5UVyAHDwViSgalYJdrZfqGlyJK0SjRE3UqkRaMSC
dtBciE27dL3hyyLlDZcDht/PEE+FqfqlrpeGqgghxB0sJ7cX+Hxh2UVU26hVANO/q2UiMo01Q6gV
ZsxpM99R0lQtECtgjuKsA6MOoXGGH5V4rzPXUaL5qOxQ51ce9er+S9NZG1L96Npg4DJ+MNJPQR5N
lcvAhCbGMwhBOWZ4aDTb8zijrE6VUSKISOs+FMVRPFoBFE4LCVb1CFoA24NjVl42zEyJ7HrKFlmd
X8KB5icHOS+bkikfatIfBw27waghr6G0IWY9NQa4ZXPJLvERMoDESw1iuohGtvmePJ+dBr10PV75
b4sShklrLF0oogEgtvAH7fhoa17xvEK3qZQGi7ScMzqtzdYRddrBLjZO+i5LPYBG2IF6tpJ7JNIv
N36mGBBGiOrE4QWk1wPOWyF6EUh0LAoaBYgJjXByvzIdOwC50GZEKyxyY6R0Tej+GFPpgZKj8xT+
txJrGLnzh1GLGH0V7ox8ax7GuvY2L2kUBqcDth9G4NEQve6yieP6Om8nu4TcFHy6uDjGDNGa9vop
VUgtNmC69RWzzA/r8h1FVrgOOscCveD/Pg70sLGLewjtDO+6dY3RqpaxE5CsLF/DjzjvYzFP2h0n
Pc4E1Qzmv25xHllN8QrS0dRqs2JLK5mX7nrr+MUM5U0ZuinAnYkmGU2R00d4+F4nYIYM6CL3d3ch
GWYwfQnJA4MJLq5s1R62zHEBAbCCaiXR9BRw+LRAN4GogYlnI6HAnRZUFnrdEoAgbG5UiJBxLuc4
EfSKEuDu66hzt5nSIOv1GoN+dMxmv1EyTYBAEevywL/FREXU+catohj2bk9y81Cszp1gE+APJ49a
bL8hJY1LUZWUALxr71TlxcWSDkgq9sjyKs4y50StNcgwVvORPF3Rdq7GZZyjCbVOBXPEtWAVn6JP
ydZywUAuEekuaZrCv+MjuLBXC7n4IytoAcT63g7TE8FxjoetLKvE3cJJUfJdLd/OJbYO8xJgbWCs
2RlFabwD/VKICGJieiJG3JYETV2Rhl4uA5ex+tSPLgdMURJ28LpM6TxaAURyCFBHwFKzKmiGyPVH
ZIygPhm/BshYpEBW+FzPz+2oth+8+Pq+73G01TshAx9VqwrPO2aaosFO7P+jh8pcVoNkHWXY6F7H
y+8C3SCUWuN67fAlxgwyWFBOWFeu3B4td5YfqjSEhsAsM/zX3ZEjOB2bKdXjSDy69GC1344VHmbi
hbp8pGq8Zx75gZpWjj35aJPiLqjHm2Tqa9BokvlIOyzsvpoxgkI9n5rwY9NUF+yInCmo4CwWd+sb
GqA9lDZ8em2Xe+NtXMbKN36K6e125kmnARVw074jo6wifNej3qHK7kNuXvIgx7pvD063kxt5vTb0
1SkwQuOlxCWO4mHlPamRrxFPuKjvE8V45+SM32ax/SZr9s6fOU52V3rV4HREjsO0LuS2iecg7M34
idMRn+F5cyLuHeGFa5uAtjx8WzdZTMfA8JALvo4/5VemGpgK0mtZ3M4fnQMcZEwdqmkvj6LoPnP0
9eHbW19efXtekNrTbdhYPfLmKLoIWBpC85VxMLx+VpnFCQdGwVyOANcK9A608QlL4Up+3T4Oay7P
6ZSosrR1knyR2cUhJ+1/5kTE0TtLdoN/rAv7vSAHLFFUomeKgN5Gb9qpB6pm4oopVubDFv0K27Oo
RTDmq2GLJRuNjz9XhaEHmj6e4hKOHtCYx2G6BgVcZQEIRF1qNkg4dF50b8uv7LDEjOHeJen9PS58
pMR5PcAsLFi2wYmOuxMMN4pUUycRELV+zHp0XgNOEqchr+ucrHTzdS3wOOAisUdPbXp9khjhlVLi
bqJTo6h8EkaDu+F/HVC0Ys6L5C1i2SWyXIJ3whqQa6RcPhVK6BQlUkuR/uqC5UYvT5WO2Zkn1wO7
1cUIwaTGot9TOw5e2doVun1tMa0XdRoHy+bRAaEyJo6K36tb/K3ogO5bTQJn37OUVSPYpGJw/4IS
h1hOiNrAL2VVyudbrCxb3iMT9OdR8upclZ0Qtu+AYMqWsbGUOUir+HjkJ2UK6QI7p3X72ruAbGwm
n9nTzuS7/YCwCrXy2L3lfhjH65dkV7no/KnvWJtMWDScDAN8PJ/BffpZmxA/QymLksh2cwjTJTqC
47v9dH95fI+UliSivN5a7h8VOQnQ0RmxiOmquSFodeklR+yGcxOEiv5zL/8DL3i9rIH5X/Mqqlza
v/keCoAR7BiBp0xLInkol4ZP0ZajmecqqUFb3nnxBlG9FDWWOBHk9b4HAfcz4xE/TnAoV+LDCSPg
H7KiMlxCd3x/vHufICDHC3IEa9nKWvr7Yf8hvburl/X8SkJGTAbePU7eKkfr5U2MQppwcNQE+vCj
S0VK6ux7Z+qN1pekxIeAlMxuw5JqCv0s/uNj6kQ3rcC5BxPK3fe+ofx+EHHNsODfSjUAYw7S2iBn
wM8LOXCG4PGcglWW3XI4Rkkrg6o8/PJ9sZYeTshAWDMdpi+SrYnJGT6ZEa1Pfs8QYE/ClZCBHrmQ
X2em3f+9Hl2lVnPZVAaZea8hpUJirjsSmiigLAM0aXSXQOURppo/8/iHb/6WkSZhE8r1av+ZcpAW
1lWGiJvvg7Xb8JBWqAMAdxdSlv1wHIoopJ/oAfqwvXFwl7DMPV/cd3C6gQ+ADRVYcYsJvP349xe1
hSYZfU2hNE4toJd+Dpeu/FzKYYlNFLc44aU5/YzD1XIntMdBAZcFMDW4rYTruGSO63a2aJRFGrIK
zBogNcPBqfHL4Y7PMT7/hmmNNn7SNXta99aZIhcR8xJ9Jmv9mxDYMf70mTsPmiO09IFIf96w+hdS
vOfhi+bRPCRXpH2oDgg8do3xjyOl7xyr4JL/zG6FNOjni106UphMvQH2is/jIZ7hoCOmj3SNquWr
gxqsqsexhoEfy7MX7TxwiHazgyFc95P5fD/uoyKNW8NIOxbmr1VTBSeoBBpdBZHCB/ru1QK3BQaD
wyDl9YsWzTHjy364RTnoMTwvPuvpfN+fYoNcWZ0cgnjtZAIKGmLTvKRQIIm1uAy9P5jp49d7qk4a
g2yVIb6Fo8poRLUL4Q8LxSdMHeiZ5PTPfDBRbq8IyqIKPLXLU5toAHbXogH7FwKM22ORUdaHki4h
jhrCyHOasNkWcZdGiy9LqQjVOXBQCikXKRUkHcBP2Gjt6FtpdPTueotB6eH1RH6kOgb3U5FOWSo5
BDBQN5C3lRNdAz06MPU5dRYKbTCsUD5S+ieCkt4spS52yz2E6A3DvcSGbE5MKerAdCrw/C3Xr+nQ
SdnVSW/+8uOxEoeFzNch3/gWmSpycWnbmz+iZVxHnvxCoYrOMhvJOLuv+k+ZYCSYFpYnrlchKEmp
HfXNU+6imgpgL3ZQ+eC3D56i4Qs/Joa4AZYjZcDDdpAVvPiZjnMw8PiTbb4SAlatCG/njDrk+Vai
7t3ACPG/eCEupH4fOGu2iqPZ7khzd2KkcySiNf19XV8AEftUv91e5Y7/A5qbGsqpPGILHPXnGZp9
0VGti5IlTpLYR0MRjIzzAYrKT5KlFMoNCbX3L+LByJ4Ypob0GqumsDTZCGv8vOYIfQi17nYjrJ43
OX8hneU5FXN45hhSTnLRAuH6DIFYHLmK8FCwLrDTNwBuYkP2oYiJEhAKGyF/OzTlc+khCuP65AUs
J/1qlZRX2TY8A20sh2hux5IrOgLItxHfBDXw/aDehPVU6hZy8PgPKrtg7xTVST2H5RVlJb4P3Zfw
9EbhL1f+LwMDhdmApH+6Ch1ziTDuVhiD/4M623g4Uj8+Vmb322SUvWp96LrPklUzFQYjO+BPejKn
TXv9alqHu+AWnHNbhiP+ICdmj3GmvAH5V02x3G47PphWQUI10NiefoCyXBfLV9PS1c6nozWwTfEa
Rewl4CJTp01aWBxuAr00tA8uA3oyrBTdUMDXWyKH0bB2b/+ChF59WlI7VunLoRPDzGJ3Czymzwvr
s/2UJusKxPCDCbyITXkc4YgoISf1svuA/RSJyKfz4C1Ya/q5KnnjwApfiJ0FE3bQXeZq0TgQTYjR
hZXO0xtku1g1Wkm6SD9ZUvHJQI7jg5QL9D2PIuYlsVuNtbFYH2wTd2UT5i2R05dHhYl65GXAdIIp
ZAQ2rdG3PMkFf7ZEon9ornM02Aux/ZCjl7L2UhRK1DUryDs79kQmwtbITYo5oPUTx/OjngIoM9+0
RaLOhn1FxY5m1OyGyWztVtr8o2evWqykw7azd7RFG++Pc4y9tqzRmLQZa6nRbpUDK++rILa7qsaJ
ujsxYyw30sP4z9tsFEzXW1f6/PRBdAsDjSMZYPi/Nr8sjimsWu8dS71oYQIsEh7RQp9xZCeQY/Rq
gXn1NWNfP9vnpV1x0A/ojs3H7iPbnB9vMKiWP3ts9CuahbfcxvRoOPtkazgv4SpWbwXMlxRrd12h
9WDksZzzngNUvw+pm1j6GD5I9yFiBBvdFczEEBYVgpmX4BDpsmv7fI7Rvn22gT2BC94jN8J8V0pD
I0N3FQEypPcDHmizDO9ywd3iC3ohcSwdLy/N9kdsiorfbSqLJKO5FTAknh6bJb777IHrTgfUG750
I/YYKMcYnA7ZUEdQt5SybZrjG0ldNEOiqQRK7rmTixFsqTia7z2pfM//nzp2YMV7bnh6FYxfNK16
Eh/FPQNUHn3ya2EsjOrUIfExshDNX2jSMsUy2iaBb7dL8H9Wt/EPMW4Nn3/c3wHibPewTxxOLFod
9wnSatjy86j07L4lZphnm0RaIDQTF7cVTcVfV1c4M0JdguTmOw9Gqdsf2deteuPivlQn6B+1OOwz
z1EbYB04wmTVzds38lEWl21Tc0hHQmBeUX2AoFWD468sXaOAaVqtnpLU6ZC8bW25xBODfhcIawc3
6a32blcYSTfrvc0ZB5x/cUyEWAWA6FyR7Au98MQtAy9Cu3ODkG+8PtAU5vIrciS0D8HzU7vFPLt9
eLamuFGEyllINLF7LymMm5zmc4vseyrUSvCxCTYcfKjNRHz/P11EaVreJqZ9YEa3044L82GnvJMN
eB/N8aBXZBI9QiuVViyRMxy91Ihhae2uUrxoYtCzTV4ujkIKDOE9HuNhshqZAEzSrJd3OY7h5UlV
T3ujNmmMwB/4MoWLBpMjAijcagqpYiiRQ6len/MITGyg6fsy8tQQ+TJUBIMseVWL+qaFPCeW2eZf
YhPNLewdJvia7M4+2tnjCnWTt0+QlLTzfhmS/U5QSKiQKP18ALnzrXl63OzRS9oVke3OWWcG08Kf
qUTiGwqjeLwBDi5iO2r7SSI2ZmnRlPuOgmAFiqJI58dJNwcj63AJsJh8I0HHmqTHf5Lxj1I1RIlr
D+4SluIBqM4ZYEbpoUCJDXKf4ax2CgqSpldvfxznbje7NZd+V/NKaHSaayzioM4hfQ5YC2VNPdvY
b+guGxl7f78+pyIkaZCES+xSaUbyoeybvY5TUXhH7Pvr70nnP8mQXu3iWHtlAXEH3SCdoAkHf9Tm
w0jbFlZjM+kutE024NgU6lfkKeVbqR+CKs5Nkgjtbd5xA+eoJyqrMDLzclLpSlvt7G1OfA6948DA
dFH4AKeFbALKElS+sKy/JZINZJkN0I78HJrjg5rcCjb3nOh3QYTT+5gDZSUf5UKLXOa6swx3XRt4
I2NjRJx8tDfxeOSzOYITsIsSfJaKsG5bjEcIhvJGr8Wlso+c6IEBwQAJaS6O8OytozRaYhr9yEDG
mRI1KBpbOyDazO85Hs6dwpMuMCtBy+sPrkgnl1gpKDtCwnbGTEppAnMgzLK4Ao8QaaCmGXQtswWm
nUIiyqgMt4ezfAjw5kw4eb5nL21gv05hSxQK7Hj5Is0aZMZPqkxKNO+FuF5m0tTNlt2jcR3zkmux
WA8gk3wgsBz95SuYEfGmPOnNrwatVcsmexB38ObBusZMrt6euW/z++IJYhL3/h+ooGD2oQX5lpoc
xC94qlZgGbIEwBOUjlhG3lSTmsm3G5OB905CjyPb2RAnUkXusM63pcUPNqokn4NNc3GWYF/mT9wH
K252gxBy5UoYiBMm4ZseLDuCcxB0BfKNbm0aXX1qyhGi04RICqUgmqYhANfDMeHLGyu/Wl6Y2Xrq
iVWZiRsUDaDjmrPSOlNYgg5G/a38mUSCeUZYJURG0zX6MuAjnwn3hd02ZoIfaAf2YwvN5Xkc6c3G
Pf0N6p8MiixI2SQ+9OUqqRbx2D9zNzWseXfml72dpmKxnm88g+r2vNc1zGlYnyQunv/E5z2Vf/el
mJHcFctSXDIxy1AAXZm6AczQMGApXgeB0UacLrNF7YdUq0/0LKGk80AZ40TyNgV9aTQC/jC/1sPn
2nvScuHzofx2mzG9E3ZsmEbLDNZNQjrF7cRboXnrOHuWBZtz/jzWQ9G8fYUeMwVM+bp+mNEkrA0q
TbsfjDaRW5MHbzRTzjNepFfczqlEoscmt4eaDf+h6239MQ6M3axuRX0aaeleCKjUlM7i+TvS9W8o
GEknE7OUoyUKyO2Z1zBDAufkdCq2zLcLuXri4XbhuMaSe/ubQ1hFIPqie92cEWgzpQ3Z24gaQ33E
1u6JTMBNHciI7z4GW+OVW3XZKp2YkAdeWgOUrnSzztk+CM9v8z0B7XPzPaF+814Jo2UzssJF3Lsd
63Onmw8W0AgBgWwW9OK48N+CvK8eiGw+DCLipf0cjaVqWHxMr2qlo2fsBmacI8HbErr5o/njgzUL
G444AzUANtvYPV5pR3xNeSKKWp0kYbpG8ipq3UsuGZDIUo7Eyvyr2oF0Mdp4EKDEQfHdnUs9zovC
nqnxdeN4AC8Fb7wL3hx1ie0CtSYXn03GOhmXwO7PvomZ7tWPHyUyJgmuvmuf2n4oHtRYw4RaPRa0
cYBt0Y1zZuFRjlVN/0kmnHR3xwu6Z6ERFiIvCvVnFdPXcGGvTsP89e6VQQEL2P5VQsqQMClqrDXb
HlbFfMjLSPy088t2R2rc3+leG/oWquXfRQ0gi6NknQMdUQJYVPYnup/SZ0I8OLqmGMm9co0PufGj
QuVwJiIy7P+J5iWDB+M/3acdW4lGmDj3TA9r08S3gk0NuH0JaSFQunclx8+bdRbM2He6BQKLjurr
YO3bQeARZSjxCfgTs7x2HSs1CfegOULvjOV7VmltXOW+2hCc/qYA1Pe37PkZz3U6XDHWkNFlUfzd
GZlRqIXQWvapCxhpVGBUi8M7ZCmtO52pod8xtfBmAsGjIqgyjmULRoYRVrL+TWJFGWJO5jqxP8vL
6cQCcnU0KMKzrSRkI9OB6L/O06/mvXt7ptRwXvH/hIRQdFXqEHZ8pkxKE5UmL5sePz03ib4L7nGI
dPrK7qk9n5YiE6XTDHwYlORnDI8AUcaJOZ/vA3sV2H6iyigcYKM7U+HTkjsZ8FGupEfJ/8sek/wo
WD+h5/3K53cvV+kNvXuZF0pYV3AF63hJL7bmoj01iw5M2XADlZDsJtu8Iu2W1O/lNOaW9o8dNh7x
f8h38nWotyp9FdgyKNSz/iFM62v9YDae38KfVOgZwwNuMosRpd+oxs4OpNf9yGkiaFSe0DvRVCeR
M033fCIn86Te7RQ11ZRIdWxTEy/QQzEVovon6rOw3pRdo9sdI+IcJVsGAfci8pKLFaRduBQaP0MA
ievRkhKqUXYKpyE8gReQ2KWou2RAEFtz5Z8ZCz8PKdBrdL7YXqiEvHSh4hgtXY7VW1lm8rYwliph
JalR1e9ahWyaamLbBGIovMQ0i/d/jfgT6cDAkWfkCQEuoGWr41vn2Elq/4O8qKmSuMTkPvjQWOAH
XspTjDZ+KoCpNRjpVYJauUH2C/BKQF3odbIzCZ9oab0SqjHhBxCXnQ16kYQGR1+iGm/VRQjYv8ib
DdPxhH9I5Wz1w1hICF45ja/4ETerB3oxnNcbXMnIwVGP5vo6XiP6wiOFi9cecLDsK0FB/q2p2GCC
CM2da596QOjyLPJq6kHoGCwTdRV/QhzcFyYIvxOnRpA+ewSoQlvko4tIAYbkksgSgPCuDzjFkb+Q
PNXPA/EvERVziZ6R6rrnaLMfoIAJZByRVhLofFEMggmGxxFZCqM7B0R6utbKUwLrsblwtfYtjICY
jnO2wMHF6lV2N1ImJXsRiMQSAOBrtxKKH74AMvnHHWnWduboc+6d01LGvueDKkFperenYh+fOubq
/7sEL6iI12Yyne1801neRUdkstUUl4nfgE66KRZlI/3z79NW3rG1TVLVWhzKoTC9DQr+pGbHSSmd
ZBi6Jy7Vm7ZrTqlY/1eXriAKOUfvDw2uBBCFmc3mei+xG1zRXVxDEClJ5kDtXpSCWktvI3Cy+y6s
1Pk5K6cLMpLy7XJKtoeOFxoh+ddAbh/WFiTQK3FMgCZUTHS95q5EDGpgt5CrOIXJVXvYkJyI56Af
j4wz2OXm8c3HWTtXBj6lNiCoE9WiKElftmOZoZQN4iDOi3v5cGCAWAo7WQbtO44OE2I9gvLYltTR
fjhGtXBMxtPyDqSbXVN4NsAExudKG0HfIfgssrIOUKCjCVD7/BTQevDG5xX97M89KU6CxxAHhtdK
13ghALq3vvZ7R/9kLvgB0U59IWSAmbQ/91P6hoeieDoCqVM+5N3DHKv/ubsz3gPo9XuEHreI+qRh
V1CuMadryyZdfWiL1Oom8uLxZcXzu+ViuVQPG7gsNnuVupC0Eg86x+vIii2CectyXYRR62yxINo8
TYEpSLBq6pqFk7/d4UNbhX8E88nCunJ/ImAPnyRFr3s3mE1XACcvRIDSGBpqHqAmZ4SsmJdBEaxN
ebZqNW2JPmn6ksgnOvPaeuMgh1xtcGvgv7FKuN+Ux6mtz4yHGYGItmu6nTgn1YN6uM/h0G4xoP12
mP46J9uXNioAyggGEMfLOwkMtcCz0sFyOsMbJAX5f1pJQYV2AGYI6fpv9qJXm2OAoBvX+3VqlOrG
BziOYA6Kp1efZfI0OP9/g541MWgSSZrfKEd5nTm4p2mNjW0lqZaI3XCUx+u00CpE+O/B/6W/YEB1
gApxE6BPHptLtV4ZrWiWYu0RgdYdCVTy6cM8zPTI02U1A9BH3Q9sPwmvM++59gcajYjT8mRFMDcj
YDuVSn6qIDpyARh58AnGr20v9uvMp9I7kfNFY4qZMMvPtmZv/5k+pdGvmp7CseEx5vTICzCmiLFS
Q99Eezmp0pnK1Qe/MDm2tFGFht86yq4dxdEBJP5HjdfHZ5mNxNENsdxLZAbJpyER+my7M9RxTbhf
0HGGYCpkbTxJey+6Uv6O/xRi4dh52l28FsVCVpGpfJXk64cDti5vTLfQOFdQsSDK5xo3e7gdmmCx
iNSwM8GuHLiwpVh41V0PmEZJZonGv3ucRLNn2o4QhlJ5QYvFTFeL92hzYqk2KcBETrCgBBtOY+LC
T3MG3sKs6EsCjlDzLOLHefZ5DUac4xxAFgzUEKZGakI9CRANkrmRtiJdmuM9b+HKFBK/nAG//XZT
O68f9Ci45mzeEwHPoCksOAW/2SJjP49VHHxPZkXim7PQXuI/8gbCfUPEsfK/PViDDyxGPOgcpM1D
mnFPAAL8w/kpm8tuUIyJ3DkFqHX4bSnoBXJAzuKXV+AujQR0F1Pr5f7abmvffIfqrltmOcEH2GKO
LXSRQuON7+r/+FMFp93AAi9A8JAfWoxUq9CjM0wM/SOZWBJm6g634ivFwsDK47QyfB7n8ks2WfgM
7LjHZrH4oUbbIAPGWYfnxmekPABeHJZ50/X5r0jgaEOAXmqB9Z2jbD38fPD4WD/J3e1Ycl9a0iRY
bKYg09fJw4hN0mmq2w0ui2xvSm7t2bIIrD2CHE5M9QekB+4kVZYLia9WdJkX8wss7BO3wFpIOPFs
ZOaY/qO8r5oeRJezczJ084rNXZ5Y/NFx8/ca7plivM72WEC8sLZu5J8/F4rl+uEIheB05uNmOK2a
5wkxe3SILa7nhxp89bfzZYKhQHu/TfL5gTroYQXwCNDAQXrpJw7dcY7EuwfzgUHVxbS+cy6v4oXO
BzajvLt5btMrAUg/tXcVDAvzZnHiWDj0WL4ewknlvI46Xap4mfX5JjBYfNWEGNjQEmaEcFV2lv+H
QqOA7T6hdtVgg4+7VSN71KK7IzSrGS1Irpi78yyJ4EdehnlKItGBYwWJENZpuM4S3o9fhRq8dcuy
hdyAxpjzW28xpBV3XCN5qlVGx/7RY5Rnyp8bduvprOtilM5w5JQmhBoqKDVwTWrPxIMpcarZVAb8
jQmnDNKV+f8lyWgylcZBckM2nyj2/CxQ947vZzUjoqtWyJv06o2mf5jzYPLS+MJplHXZqfnrPzhz
UnbwD0aZMvVygjFVGunp9Mlz4dYQ/D8hgHVVrpi9cE842kN0Hr0+IgNCtK4nIKl1Dfu6+zSIvuYP
xfdbBorm8gvcUNV8iZ/o2WvUy3W2RKsDHOTQZ3i7PmPfDbChMDAu33kyy+9pVx9iq1G42aHKkjeL
9tjyrYjVfg2xr1kesePLZ6IK8hAyLXT1CcrCSTNgQvijofiAFfFzUFTg7KsHLuqN0En8DWM8K/F1
SFNoErndqMNObrIkU9Tz2xiQJC+UfEU5nZqNXIr9TqGyYTG1M3cx/9Y13LctvbwfCS+Prf2aTRmm
0fGDeRS8OW+p9ZcGXEd+Oz1y4235XPoOmCct6uGdK+b48HEOsHvQeSk8Y8/TezXJinuRNvDYsp2T
sTXpt83llr0rtAnJ8qK0c6pIaWlYN8mhNGQIo6FCNPTuYiWNFqPwdYF1ckiBHNGzqDZ6nY2X2J3y
Rf2I3wHHl+ax1tKWBpzCtoUfvLkwn4qgwjJSyYyuaSpYgv4qv3kwZJOh4bMAZcUNwK4fEJL2bgly
0//10K1HqVOb/TlIeO/mbEUhw87pSRQv/32X77bi+7U+gtXX5E0LGUsCTLdJdmsErhf/TWt+08bU
LOEHcl2C55uxY1k2U3R/xLN7q5MABNhcsQ7138XTC0DoRFZwidWkGD4s6ZwNA0eq6UOQ7hmFANMh
ChVaSgtzi2yOAR0cvt5Jl2szfsCb6hU2ul8xNESVdiytn842N2iL/rB/7pI44QlOEuSGGkHqQj8d
x0Q3uQpKERTNHhXWPXAplTcRXLIRMfBpUwx5oDXx+H16Bh8QB+lw7ubkfDD2diSVPA6dxrHxynB8
3BYx9Xy08ZqJA8f478CVa8jliVY3LTP3nYK5j/YvEQdacAKUCAv43j4exL5LM//xusJYWpYQspuG
oi0EsuZ2B87LYWHGqnFJb/y1E8fchuoiiN0YYtAvHFPpGz8Vn1k40OuDKmI9Aa897AKWyzoee482
wb+igkYbGMo6LKc/AxhDemYojj0FwVAN/3Fz8MdpDKRSqk39OplfMN/uh48PfFalVTN22Djbn0MM
fYigsShK7fXufupqSwQ3S9Bi7Tae3L5j71qtEx0C8u+qu0j88JJv4O6AJj7kGfHfq468hMfWtn8c
hJJWrg5qiikwbefdfrJPa/mRRbZvadpetGA5fVxuOpIyV8SIlaVKzHQtWUacANuZYpcLpmBYOgvO
b3ZAiG4fx7PB6uRM6wM3W6Zr5xAv3UuPYu+evxLCB1MHfCDV4MYmRPnoKE73DxSJjoomXYGBS9kb
PqohDWvvgj91RBWkKK2D2wYlmRLMotUes+/O1SJfE5mG18xwq4lgx9UbZ4DkAn6ax9ECpfRNpC4p
yb6LBROZHZl8XoYOisMZkOLy8d+uN0qN/1tI8syEvQ6ZTAGa1ThoZB84kb2H56tK8UmtaYYmOE1v
OdrBmCY4EqAbbjH8v+GPLbrjoQp+VkdS4Rz7uJgTdsXPOXOFLojgjVoJeXh3fj75E77r+bLJ1vZH
oR8TTfZC/750Lgd6GONRw6PjLlyredJ2qBZjjA2MfRMeEmwC6rXitYwww/40whKQ6MTTWMbppegt
ADBA7VWX4Q1kAncJyUw9PevntP08v6fnKb4A861nhpcW1KtkJAZ2g3vjIDQXfi2Bvit3pkPopX3S
9f0RAEJW0eA902nyJ4RMoO8ZrBiayzpByO8m1BBfuCzGbcIQDwefFpwmzF24Yl06PjoJIoZPFacv
cd4ATOunOOIRRX62zXSIY+rIcHbIoEz8pevHbdU5n/oi2pMadnRtIueIbXHvfdtIKT+eXjcMdMgy
Y91ROxxL1mA6YhiIun13HmmGYFgIzSheUKF61ppx4HjAF50MdAa4velyy8OR4I2Odqv+fR8up13V
1+eMxFi9X35k9EFivnYOXLRaP4VjM113b62Ry4Jy36/3O0maS7Ic0xyFtBA6xnHK7s+o+AuitR2J
hD4U+JnKcYulnPwPMRAh9kbCtI6OF20k4A63ahtftBEOaUl/3IQbuNXk2dm1iQAf/LAd7HL4oL2J
MNqYokOrRH1+IA1dEkP8LXo+w4ZFmQqfRSvKikxjJufzIYIWrTGmlzLx4eJDMfhEsnlKsurwfNuf
B9DAQbll6WGFkgBwGj3m9dJU+ISY3PHGlGb2uyrCKaJ05DXpP4o1GYuqig/4i7hJLLFZFOyYRzQK
h2DGnj1bYl526vTXaZFZNTFCRzAzvP481HDUYE+xN3rnOmYutuJZuCvTLLABoR7eWk9Eiy0l6WZ8
pZl3PXFN2QQPp2rjXlvSWInhGeI+X7Kma1URY60s5hCyykUdv0+EIfhPmOtkm7nwOlOQkt3lb0iY
0Hv/2wR2DeL7NDY0CorMUD2b8hAt1F+Q5Y/SzE8DSwGMturd9DLddggu1eb2CSSklTs8kGisy1Rz
N0dJCobKRt4EoU6Pc2jcmCEvWeGUuq3NLc19pAC9qC2Vv/hbwmUpCmRvHYqN+mU4G9blfgUWpSOr
mOcgZP0KPRAusWrW5FNcJ9vhDUAEN6b6wLaqj63SzJ0B7fTAyJpuzSgWGjY0SzJEkgPPqoAdRgbi
pudILTVAJ0eeCz5DPKbdLr09Ia2ccuMMp/+crYgITpw2Gcoj2S7d/8WFt5JtjT8xHvhYElvkDHf7
7XIwZoZrUJ3SXGJee5yEA2vEUHsSOCTT9P7IU3coQQUS/nmEp1d6C5xnTPpJfym+E/Z4PgODe5ri
cEhhzRS0jdd7EZdgJ23ZK98ELG9LQ6aidQBZJDFb9pSJWYNFzKooWbb/k8J77xb70c3SPEiVFKJV
/JTYjuGvOGuBI3aTK2LT2ObiLDFJH0PZJaEFgPNgEtmd+/JKqxAUVV5eQEFg356JKEz7V1jqimS8
A8R1fNlFo9AmrTXirkKi2JIb0Df+HbL8D4vn1u4t4CcQYxIqy5BJljYgCPi2JrMaAJmpT/cd/3U/
BrMzqvlXffvwGl8N80g6iGRyH6AwqUug5K1OrviUghoCHno9L7Xxlz5mYD1+0tdst+Y4elUyMRmS
k+k0CgTzy7eb4SFn5393FLArhtwSqvYPE9dvV5Nhrj4z/Bqts78Z0sK4Hi0wXcqFUvFbZALyhxWO
/zpOmcL9azfzx5SciHHvotivtLgXxGj3C5I1E2aTZnpi5lOBXPulMFf6gpVQkTwHY0soG24uwxSm
s/bBFiOMgrTMAf4JbMDkD5jGlCaADNmgBJF6h4j9oQTABWj+jcKsM2uaGHC1NBBRDbvVm30cWCgs
YoHvX1SiRsukwgqGHFGvKqCdfdlsLJKWUreTkgxMe+zLPpDYxN5jEIcPJe0V3V/RfX4G9JBCeN6B
8PXKwnEg9pSnrBUlt+QQfj6U1MN2gbqwO+wPg7FJMQ6XNYpGbsZY2LsU4brJlwYcKrK5jJWIHMy6
9dBDM38sL0nu7F+8hIViKNpJnXc79r7X/AKz64ACM8fBhQ9rthZ4oCyfvDzbtbZlMx/wyzGmH7vW
4z1M+IdhZE7pmI2BHtyzwJzvuO07v8Tr/1W+gaedmceQgdDQI1pMJSJfMgqh7I2o43bD3R1hbvqv
qSjzEdcVD/qcZZAo58eL03Sf38nRWchW6eHBQrGfWaSwMkY5lA3CjwRwTurzCFld8ytx2L0CzTHz
ljqz59RKrGwdjcO6dQK2UIuyHS/p2YtZJcrh6VmjXjp/zjKGxDVl77IyI01E0YEvH1fJQKM+iJ4W
qc2XIZ20fOzXeQxJk4LoM3f3S9WzrDz0moSPLkcX/Pr7d1ssO7i8ELOPFyzOp2QKlKaLzWci6rnf
TXN3o8TmvtGRskRPhSIgLreCMgSpuQcM5PBzKNWxWjEIGJSvwHfJMsEvm/dakYlHr6nD7zmdBHeL
/Q/2g395mi2zT67UKvJjraPBLqkqjQYWVeHYAcV3QLwjv35xfxbhcjeiLDvFC+xffHHa6AR+KrVh
DDQsxzphhDx29W3u37cWLo7pSV1i4fhOu5W5pinaCYuB3CFNZktZvMB9nyDxifNi54nDB5LWGNeI
R0cFskuJOoe+hEdIYFWLlaFKWuIw/HuvCghMYSDzLS0t49jCukfjO7g4CAk2Qfkyp/axvAx38JSe
RXojGkuQfID6d1pc38Gf+HvGIBz4nlT+h2FFEtqJGdpUaX0kK81tWKNBOBw2zTi/TYIX4qbyk6vL
lvvqlZHo/Sw302VkrXEM6c++GkgGV+GuQt1X3fLVApTv6c5pp029BH2y7jnKoH+U0CqjwiEcW9zn
S4hA6h7SNtiMTrANyfc8EIXJw3vTgQzaDpfdW3EaI9JAo0/9GWK3YiZqkCulJNSyNZt/ABjbyTj9
dNqrFBoDJ4ua069U8GrxsMAcec1GPLfzuosIYOyyIx5vmxio9siVwSvwYSj8pW2yQ6asmeXK6Nx0
MvOdfFtczllMoZ9yFNczl2mRkJXn46YbUqOOubcsu25JoAXkA9BOkEW2cM9KQF85dqAGWOgAZZAf
ISIWYoGQ181xn/mo2YF97565GJxsI+Stv4or+kS/P5H8HJZvGmPUuvJP/IF/z1Sv82+h5mPGJc7u
H4tBIPHvtAdSTGmse+ZFBFGXdvHmrbu+mP6RRH85DKydWKF5bkQkuB3zxxsek+6ZeWM7EGtpPTli
9BfqX5BUWYP3UpcsYEtCG+M9M9/mrOqyN3BEbd8C8Z9cTmvZ8ncL2gQOzfzMSzDFZWcj8ydvYWhS
+z5OwQlqypLfPtzHCz1vf3BZpD747fLEmEHhbAQGvWElTa4TvXySQZZQTs55MynrAMnXjmiC5Z1r
m43uKs8Ad+Gm5OgrR4gI6vrJqGU58CPgxcLQJvzkYXPXotE6lm7ben0BeWiR0k1HzU7Ud3q+Gsc5
a8b7ejn8ZfdRnVIGd3HNvaDXQBfirmLk1CBGSeebWdoz/EpudUyW55qQzUZVBeQbbqdhAQzcJuV/
asZjSC4I5kDghfS/fR2TDaC4uGs7n5tsaPI8fCorEgsUnoZCPcCTfoYT8yCBHEs1cFguN79GCbGR
F9rpbgImPSfob/Goq3qPdFH4OrL6kWNlymBis3Y90Q1i4DZ4R5mnv77dn+Y4R+OoO2QoKs+bsCwx
qg3ezmJiFq1Y4oNGsTKqL7/XwieyNLlf8WhShomxJfhxzkHgpT/kron49cJqzyHq2W6HZ350m+OE
LbcGvNrncDe4NKKUzpNuFZ1cQ+jc5Zx/wkKrlz2O/xVxo5g5xUdlGvDZqUfTFczG/TxRsQCshF7r
TNFW1Ad3aYy1W3Hn9a4fkMY/op2ycsZHH6LVntf6uB0fDU6TD1T7lv9fYdQa3xvSIG35hKt7tWsp
zAbB+vb7zVNhZ5ZVh1VL8gd6rkoVnwt5nmcPrb3lcSj+uH+NX4MkWKHRosKl8Xcwf64eh833F62L
OP9vkM1cBZuXXsBKuIgv+ieHrJ6icW26Hub0papuOVgT9YnERiCOAMYVaVW0AgNPXWInRIZyCJoU
T1qw5L/2xJ5Y2vcvz3SJq58EEVU/a9p/uAEl06sYRHoP7bmcUW4nakEaXnovNvZedA8etcf8gVp4
LxC/JSp32ayVFa3UGQsgV2WNTLd4YCBchpKx90DP0tjhtMqfQ3JZl+ED2JB/PswKqXs5Vz4tNXSp
82jTo7WHcvOT3VyVGzipJGjPsB6KOZ9bBh0WzaBQplOuGQGHMNn11qXpG5jk2q0s7LybHF4H7s2c
PRqB3S9avxlP+FXpBVMUfkoIDS+/sKEtYmkCE94b5VzzaEJFYIDM2nU4BA66utwAk+zS0ibEMDfR
wdUi6r50ECtQwQcSHYXZ9adDMaYORAdfj/oIhe2m5jm5kwZwJbuy6K8bfBNuPw239bqUHVI2snH0
vaHInWa9w8K8Nw7rzNHKzR0rQioic2G8rj0Vtlsgr6wekwjzKeFopHbwNlQTY+3p77Lf5UvEBJdt
Zj8u51bW1wI3KUrTSVXGbNBb53/ohKjkETUTK06m7ZurLjEItPvHlRmSFl74j3bX9BoosnWzGaHJ
kF46lBNP7Hm0vUWz24UOt9C0y9Xugz4nbvTGbJhfxNvDC8foX35cYkLGGJjxopzvB3J5GOZuR/+E
9/S0VKYfdbXljXtbDOrgcA6xRhvHuc8Yca9ZbS37mnSs2/oAU1RwSLBwA5R3HzY9eGtV1TVtUGCD
ke+miEtRHP5mFuVn0HRpSeNJWwZED0ARB2z1VrMxFRn39/nL8zHjHnx4WMMoU4unp5y+lfj7QoV0
suEr56UK2dd/dHzAG3DcIQatIvf9XP6t47fnILrfsMZB22tYL7+QMC8TdRHbSfActTq67T/mTKsf
iNmdoSipXKbT/1kgnMw92O3IBYbGBSNifar6RnwRS2SjrbqSwUsvgT7LPWO6soF5u82rdlIW51lH
eVAp9VjFnb8nqNUjHq8hvM/hnJH1oqeNiYq2nYm2RAUkgO8omUOeSMBLk1nN9wnZBAblxtiZCkN0
GYSz/+HVQZI/fEoSh1vzK/xsYuPhk2QRJsPUckqvH/sYa2xzK5FoHxjPFtLymK//nvfjapjy4bea
i7f6IG2G6rgQwDZa8KETs4vOV8LUSsBFByCnO2fek6/6gt8ojx1nuqjzf7uhxgNtmdQebRT9akDh
dvGUT2MelG9EM3P2ZwSxGn7cSDvJa+MY2gN0W9od5o4GtzdLxoIav7QbJxopTiwBwqw6+keLniIq
Sqvenh9GRyKMkxcd0rpoVAPlKH2ugCIiG5zpWojOw0mBbiPF+pyL3J3C3d6LutGquIgDj1IWUyDe
h09GJ6YXECaHWQ6PNAXJk6X1RTGSq25eRsHmHAL0CJn2NUSIdWA5pPi9jwxctn081ccFyVfPLlrk
qKgXvdhkiN061z0pduJgzvl2dEvE2+u5Ufy2D4rKm6eQY+Xn/h8f+feifWgutuyZa1BQ5/pjQ328
xS8Qf+UJoTRPYxH4QANCWhh+b641Qz0vcO8iAQoX4x0KEOEK9kCXeB3LiU8tfWVoOp7cA6GzYRes
tZulGbQxYOZy1FidkL7FVs7E1RmCC8gC1hMDmmw7Sah3E8YiuXMuhGrTAKWIUiJAiVlbXHbfGQAq
456JRhZlTsGZZxX6P11oxa4PhbjpgB+q80aEL+1nFT7z65+Mb8vi3srAXmbGz2NGEfxdtehEA1F1
3piTrDOkLVksR2oL0LCJ18eCnxuFyPq9gqkjjfFeLZptK11nOrZv8m8ZvPbEBOJClQqdq4QTpttM
2idJSiG6Sdph8v6EE1mJ9vQ/1H40XAffHWfReWrqPhkc4Nf6+Nx3q9NDYKkFdLT9KfY1lxWgrPOr
xnxPXwJM9vmM6Y2Y2QFMDpIVq2W0jW9cPsIGxgvc4EIsPZIO0R+2/G/3CII+oUBhsKuqXRDiRvVN
tnUH8JbKyMFB00qw25CGyuFPJM9v7424ASoZXJepqdqSYEc5WajIo/mitrVEnK+AEezmxRLaTaO/
P2b1mCMU3XHXc8zVXN81NGf+FPl5diNFwO48mhJSgbP2NPWw2DqyQ9kuhzTeZxg38UyFBen2w0jG
u3YCs9bRJCkIYFL6LJT6RU0sWq2yDfOBP9qOvHXnllrJ6iFTXW7N6DZBEb3vfIl7Wt7P28g08Hrt
wq9+2BUCs34S352EQyhOtjq4a0Y8RdCT6jm7KsheGxHOdZvWvWk3osXFeHf+obFUKHYtLHg+HI8t
qKns/FcwyrAOnjiHhzz4BVuR7pIndAWuW0vvUiR+LtkK7cdIUmATcPRziqZmwjVarqnTJVP9nMiI
b070y779w7bO2ZUDF2R1XTbWxa6Tps9SunqIYmfGi2o1pMaaJfOKvWAH2y6E/79p0cXIWYqpX2l0
UYytcwfcQRMMYpBtGgdPPAyb1xgVsxDnVBMecRm2G0LiqLvkyVdqzdLeArU9hTFnmGTRcpj4brdv
uTwFvcnd3qGUNDvL2/5b6R7ynV9emC/YuS4PYh+Hv/kBx8TJFW9ASZcSd9CBZ7iJheon8GU4FJio
zncTPj3O+W5g3vNeh4Xj+RdPBkXohmwkQICnjFLJjfq8U5Uf66kUleqcI7ebwx3XZdWCpJbnl0KU
99+lTPigvNYL7KDigN+xVypjJbW7z7/nTdDho1BhKGxMMYicDrPZPt6WoZi4Mt20ODlzPXTGupEL
kaHvSFwGx5TTCLaE9RJNivH6gWWRDLunjbUvTxVXnGE7GkR4I2iW0Ts18VrBVXYrzWBKFb271y3w
bQB5RCNOLm6LwliBRzbGpLpRlQ5MB6Rzll0iCe+8inu4T10qjYJPXF0tSj/9DEsWHohGtTqYkkS2
7ndqsdSNqVP1319RFpCrJ3O9Qpoz7D4iPPyBkdKDYAvo0nXiFutOC6iJhujGtQuYwiImb1p5Bs3U
bINcT5SJg1kFjcDqskn8INd2cuuB+mocDy/shEasnOfj2pDG5l4YVb+18uSq+H6hLITTgWJsivS/
tICTR6tKyuPStSixNZc2YzU57crjxg/qzFC8O0uUF/NB2X3LUkJI9hj5uJgM4Oj4xWXaXBXN4gFW
61C8Txfhejs1dU15QVr89LMlFFfsis+bXiekFM05sxTH8y3B3BuYVwe5WlMrkU2qL808JPguU5In
/iT4vhHL2HSldj0d8ipP0tuTheQnUZmxMg9VdCUkLn7XknOTlW520drX7e0h9aRJZRAScpLESyXM
zOrxzLWPHDDlVb2lZJbhBhc435OMrjIsKPn3wRRRNymi5yjaOfWwpaj9x8IDyrSdEeVpoziqj4jN
g8FACoOAIzWrK0ashioLltzv/tHTZzpkAcm/g3a3SV/Xf1GKwbu1gFpQbZ0QzvI9PxLS1qRNVZKR
aPZIdpmbriRm5NShY4UF1B4s6kZvhI048HhirRCSsjizAgf7VM3UuYovPI2VB0kIMWQY9o2Vo3th
AVLt09xx7yJ7Rdn0AIjwY98qt3Z4f+N7ns4y14wxUhMZBfhe9Lo6rKp7txe6bU5bRa00fIYg789K
bXNRySy0Psh6FB5os8CxcCMM1Hsw8q/FMv+5A9EjEMlZ21JNJWADHXQvJ2d6xjA9NgO8/NKJffAu
rSf5EDU9r3mW7yMwORw9I/T0tubBJqyFCaCg2q2zmI/tPFhcGDQN7BbWyOmzdbCzvGEkNxiWy/c3
PMwIWoEVLIXGf1x6xOWlBzd+0uMmvOhf8F7X7TKfXhqhRi9kVczVFiQf4COkbslJffr3HE2yEu+i
+nU9XSsze0P04poXQ4TM1e0Y3h8cOkSmst4QHaX9pHPfsrhR4Vv5kHOacfZqJlg7UI5Ly1QZV07e
DEyu6qp/ZGZCqmFVRIpPNE2N3O+gvLFme+Ni4oaIhkSNas2a+R1FZYWJJ+nyF+UWLnQyw2BFl3q7
XodjlenS1AsYrKJrXxA/REIHnMSot9+KYl0ly60YINDXBOdyLVsJqTccSzeqWtKpn7a4tVJyLlCN
rnafhcQbV3QE5NA16MLPtECRbN5vytt0bVkuVUdH8F2HzRzRRRLmHr7pbfUs1DUR5/ISXRBerSdD
wCr3Q9FxBtK4g0JdIOrepsukkaP9pARORRA+rfuXf46ja64xjCidHejeXHQDohTmzu5oTwXu7G2n
X9jCIFZujxjmaY+kuso3mk/yYeZbPwkIVW/5qfsXtdDuKshAJIzo/2YpOjbqPgN5KL41E6ujc9eB
qxQ8l/PpPalqig9cgpfxOh0gADjljsA3sYJ5x6pwP44GlxLUbjG+NLsIt+6fEss9fIC0HmZB6ALG
fDqLrTmRxinY0TVE1Hkoj10CWR3afvyrniIjCwO/rUFXsx26uURD+G010KgtJYibJ6eM48lYSfrM
4U2YiSum8U4AY4gsnaGNGhpeyAGa/716g6cS7lpYgNVYc6yAAXj2sJNgvGHPxBgjHEhRP7xD2Mnw
mjv5WBVQ/w9Z+3dHLPf5qd7HNEJhdTj/By5ao31sQ71zbMGRGflOrXu9J6xsx56XqyaR6JEkSG2A
Mq8DARuWBkkf5bnjBDj1e5SE/B8znCt9eBWCZ5DPkfzLJ5t0mYZeeTrTf8uEcTElYq8icxu4RGZL
KVfip3nleQirMafSYeLCqthyPurOitSdHtd3TV8vmKhQO/XoH7+lKSea+Sl20EODnBqH+WzzuGCd
oP0Izs3PzzAIbPKG2kcC/Sq0gCav8CaVZVugbpHjv7JKMIYIwFBKLfgjWKib/1rD9TJJqMtRjWcy
2Bny5Ub9y4wHZBC2bF4VhvxG5d5U0tFqlf2WJ2EgU1y7tGImMxAFVSzb2hSH8EkFCVTl7GDHsOLW
tHvdksvhwyAzS/JSSdLuKfUYOyBLcAHG5GgVTu0dBZB1u/LQv1+9/0rBsUxnj76tLQ3yvEP7Tv20
KX9HxFV91HBl1tiDJQhH7vE9+XGzJrXfDv/I7h6xNskvh/QGifC5xvgNnkkdRwpCE2tCPdR4CHAw
PqBMLklQF5MdFSxLD4ZnsgcSH4vq97IE74Q7oeVLipmnCo5Jm7/r/hMlvbDvzY6yoh8pglH4tcic
jarqLJKWeB7MvYeAMLxkRN0J9vxnurhXrgEqoj3UlI8oFILOQOXI8K85is+HCNZwKRi+EfjD8vgL
Kyku0Jlk01KCRzWO0c0DDemYcoJ1eGoj32st15EJOtnItD59UwEX9bcgMiZ6BI2jIvR8aUud3ktG
ZVtZbYYBnHBtcvrT1wSqj8xuNr9dtgY/dHXF1ZhGHUUKtSXOkS6N/xyJ/vYFTzYmaRXLZiv7IfN1
6wNtYwaTYEujHf9+dhS3Me6J5030YCx11qFbJfOwtvDhtZaDex1BiZloF/kH6LBt9kGdvQTgtPjI
3cWVMPqp2lc4UX5+KPyHY4lj1z7xBaaxKxc2Vf8laWSUXKZJQbhAI+TLiEDyS2j6wRCqJYR6NKCB
YgOS1SOvOU9MxsD6OVneNfjT2aM+uM5L5pVE8Am42h033X9v2KEGsnwIXUXDbfL80aDOKwBROdDo
/yr07tt02/MEv2RkkU/p+36yEML8QpDnQ1Z4cdFih9LZ6gVReY+TSm39dmLMHaORvJF7zCppQUn3
hdKX0jw60DWefMRWPs2iewY0YFoYYB7hLyCzTV3aeH5s4C03Mmz6a1pS7uLAzn9f9vSPDVOjTG6T
ry5ZFPUZidz4Hwi9JCoZOgUIFND5xHOcxgtj2k584VyDuAoe0yrf62bFjMdpRC4oQMIJFRczzN2K
0DhigCrMS3eXgSEHmT5l126WskaGdlMIBMZY9uK1TyxdRb9/dG1y3Cbfe7A3pWf1BOjZtyhMU1K2
RfLh8RoE4XZXt1Vm84I8lW5Jq8abAiEoqUyNlKmFzYMHcYdqurYsH5k8NkTbmd8Cbrj/6UyKxI0c
E0Z/GGhtlCeqa260+2FoL0m9WPxschTkmmeMBf0+BbL43iS4G3z+N+cu1/tK5fOle9HckN9AszCW
sdIiYw85x0QUxrGnkjmrNDrBRMoNePRwaGJ1Gissa++ONt4uotp1E9y4nrWeyQ7zsPyszP6mcbwW
gD0K71JOReQOcVqIz8fJEnFS6MFV1nzseswvhhnZAkOGEMwT0sVGAmar5gO3ZqEzMTQ+36us5CEL
NDpf6TABb8g7ysas2STBY4JglSzqXZjgR78vakCvius4iSZsamJxcaaQzB2Ug9FNB9Wu2N8s8XSS
vyjwMLEKmDmQmhMCSEiKbCgP1N5wKUJoZCWPtJiGokYzGy5ZAAIt59ROA2XmPv+uEGLBhs0n8qT5
o3CduJuCfnpgVd561EaaChrplqFy/jK7qaZG2tVprI6iJ4wZzyJ4jJkMsxMs5P2kKjd4Mwnvz5Io
Ga5y/D4mURKauRIi5lBdx0YNFe+v+zvXg90wFKzV0k6UTpQy8ai94opYuUI7iTSI5m2OYc1Dbnc+
hV9np16LXZpo/p9Dx/NmxbKH5Xv2hOo8LtCjuhT+ipZRcGnLHK4DyWPayJDsz53OEvSwr5OMt8nh
INRV5pM5ZBhXar7/MGm/xWt5hbrK3R9yfka6BixOmRrmEjrqHut/h3NsXsUgw6wSoKJienLOfTr/
CTOS4OBAy4JOZLL6PcuqUxjsWkYGHtE8Co4fSIsudtLNCBqGB8Y0dFb1zGoWeyq+/U9qVtaQhLYb
eriAqZdAFahFrEZBPQMa2rc2wNXpBbjduflXyJW9t3OtCLaVB0w32mTGbZRIueDX9i81I72X6V4X
OK9KuGDWpnJZSa+nkXvn6rdtUyzgYY7qegmlhIOEdfLL4aOURvHozKK+FwKgzfCvVfIJNxMPV9ID
uSWYYu5zsxOdjR3j/pkmRtAlBNPur3lTwVAqWddcJEqezCxIWNe0IZtvi3QtSKeVYN6KMFXV/6jG
6CH3RZuzLzX5tNq8aU4urmEt9EsdZTEn2a7HhK0Kk6SCuWmKz5azaiyA2L5OGogLtI4N9djxrnL8
OzCROy2oeXLOn/gd+eSQ+U4QevA28GFGLshobRkK0tOs1PZ7Vr4WWPfIy6TIXkZ0Mfa599Z29TtI
TZDBZ88jKAafeZt3QOCcwbAExbdH+NRUBNqmf8U/T+goECThjRkWHtbs8HeGPkzMWTyXOf/VD5sQ
Sz+8jtroMHf4LfQ7w6X5jjbHs5tURMzyyRueqgEDsgPqKi9PoJASz6v0gaH2ZdiCDxjqAFPx36np
hbStn+6CZOuyTosczKP3jD6VeJjcU8/3HmVYgc+5B4TDU4Xg3noJKHed7afxOviyQR4FNMcIlKU1
wOg+0JnUcDNUL7TU9LU4w/1y5b7hhhZmMWh0he29OMYrWcDVNUib5tHPz8azBD7ClcTGycM5xaI2
v95raSrSww7m/IaZXTruBQ0cx3j6GcpHSbknswqJQ5zf9lAuhLVDxfPH8jv43w71zDmjui4BZX8E
qEi/LAD0oYFIqkelownV3X3g0WKfRO8ImPfd9N9PSN+MOT5Wlyf+y7lUw1krJkmolCKKczZYqxhF
rr0evz9a46SFSVpahsFcLt8SeyZTgHMV6ppVhDSqGistMOtNRjAAJDSP2z+HkbLF29XpVpDx/ZLM
iNdFIv5RlLqDp/ACdoSoJBuqjbItjbd2mIsuPiUXD4HuVI501UwwkpmEMyfcp8/rky50gUvLkzSu
0zMlt2XVtx/tI62wKXj13fFSk1CEVKOpLQGFefWTslYgW/ILpdcMM8A/E7vRYVSUwBNNXw77qLRJ
xYxIcuypiQEYOGGB5FJe9c5XHKgcBAUzyKGkhhyQrZMFc7Bz8sz+1OmCGINFIHturxM5KZ78y4rq
h5ampO4j6CA6+DodXlQB6fypyfAj6X0QSO10kZhDayL9dYQ16fctvfp+qVhFDh0rYoUzcAeV9U5l
pzXJk3rG++qeiE7TFjID5OG7vH7RvzKkG/BFO3puhTbWyz0HswmgmqMIeUOYql4vwLk6BjmA90XX
x9xkItJzhcqfZUMMQgnpn8gHuy6YUq6YtMGhiTCChHTU+1g2cHd9RpVy3wM4op0ZDog9qxRrXxS2
HRV//XJlfLi+l2Niit8SUSc8FVSMfc8f7I+w+OrIF3kk0WVYk+Iu/k0URxRF3Y98ItzFo0srXxJ+
lvx7zrxoCsJzZi2Jxz8WQFGyOxeUOlpq7rddFE10DMTKOBtZYSx0/l3WTm0ZAnu1oqbI/Qy8OaxT
BRE5cnWUmS/kGrrMEMMQsA10PpQlCFNHW1T/7rCsD55FqlI9l3MoSGZ6AbCfEJgePyCNjtnf0K/Y
+GmWMH5CguaP7GklAVPAUP7qlGTfK6KVhp8ccTWdM6EmhvmIF1zZ4vL8pGzXHh3FDQFBWBW+qgam
Ydsv6xGGF28t+FHmwyZt54eJI8YZKEvAKZP2iBucA9vTQ7tRJ4qJz2hJ8myefz/HcGzbhd089gzT
BYqQQ4MZ/QU2mcLiF5r2GCkqnSBlEbf2Xhle2inT6Jedu3Ak0UYZHRC8qPFU6FtuSrgOM/lpHqjE
XyUAOVWSsAU8oj6BwehsbD0XejyYCAYTo0iQv/QrPdo1jSfzn4Hyr0UszDk1p+Y+sIf7EPyRFgHw
toG5Bh087vA8Rkn+2ty/1rvQ+JwimhI7PzkBlZjM/Q/hClmSLwFXdpf8JiH9ZOrATm1bTYaD1ULf
y6Cc8Y+SZs4OsneHLnMwXHvdS40QAyQXnhtTKNDyh6sW8qDVTVqlhHB4Y9NPtuQ0YvsePDZ4I45n
/9r0wq1UBmg7DERCNgTLOZPZYOnUxxnFt9QcGzaEEgfMVl3iGsrvVHe8HitL2/PsKOf7hv6Y/Opi
XYY/Nk0GqFvqhqm6ZEQ0hc9AcMdutefAVhGrc0CADM8ldv0pYlnmGQ9zk299L7k5ujkt5xC35MmH
5BhIVImLTiBr8bANg0fC9IoiZ9fxfjhZMmbbvR7CXUk/l55MKO7pNjvmmwplsaNtjNHR7mksmeZg
yV0T14JBGe2R/hSZYhru9uaJmexz9+K+p2BvlaGx56tHdrlI4cEXJt5F44Ih1Cv57fc2ZaAggv9i
dwbAU2kpGZ7EGDWHXw3vUmrjWweUhXY+V39xvryUpvzk42+UF0gp9GEmftR9UhylUTAaMIGT0Aca
J4g4jaOtVExqMWyRSp0pQg3R8gHRlgA0d48S8j2i/HG4YRj0jL3vqpTfHUEi+uTqcHU7ix/FARQS
xiEwWvMjOeP7ZNvlf4ZNsBw/EnCxj1WuOKwtTwFYEpxoIpNMe2SmkLPShkal09lUnC/GnsQ+yw/U
d3/o9YSVOInWvyacSPdEWbQiq2kQkhUoz24bCjF8yzOuoAV4bVG6XshmjUM0knNfQFiX1SuYeh3o
N0xgcEpO1MHXSQOI7JXZquVj9VCSPM8VtDoKHDl5E6C8/O4OH0wz3SLHKQkhc4b2jmyENvl0aRt4
AjQbUAtjIAm5WaKOPkm+f3IO/j4WHyLoEHIK6YcIZJ7faptoaNKLRKHHKcSyNI8h6FOY2vN3uhh/
jk6MqN/hMhlVni/0isx9tGyozvBKzWifP1pg/Cbu5dh7r5uKunaYcjzlCU/LvX3aQNZ0irxsTCO/
z/Xcq67CKEquXCTAlwadiGHDmTQ8H6bra2WeMXl18JZFVPo1rCshDWwOL2TeF2gm2uXhZBYEgbv7
vm1NdPN2lGxY9UjTdonu95591WP4PWDg/9b6/aiqmabs/LT6rT8erZwztMWdxcnVYBaTNry8WnE2
xOh0P3XTFZiDw4eVEOBR1/nAp2n6KFOKAJWk3qtT6r2HynlU7N96DfjxNe3z9/m0Od7Pk5LUGjCI
zr7FAJ93rABZm2Q7EIOpI9Zdw/i0eQ9T/hldhTycQuzlKfqW3q62Ud3m2Qi+jMI4hHqZUihFNkDs
7ATX2JbTKZWvUMSvDUlrhF496SF2UArJbo7XhwdDCSYoet+tJUTvS6E3EErGyk6MK3nfYduH7Ah4
Wtbq+iDEml1UyxzJ5Tz2QqyxV9S9R8gAkGIIm4lHSyxEhAwW8iB0KowLFQE+DiyR8sz8DdsHyf5M
NhlSlaMMvBWF2r9NueYpVLAI9VfmBmkJ8PErC6eRaHK6fP64h545SLFL7uRQzksGlzqKjfeWaXFv
D+b9NB+9mYl4yhsNdxORXmS60551hvqvpYKLbDGxGTfE3t4aUZhOJgLsbm1usbwr6BsBvEBKTsqS
xe6850mBgpblOBkpjIyi8IUmkWI7bpN9+KgB1gq+Gx7ez19ONGH7yopWTBFuoqP1j/iqqbCj3u7U
yX4BBhmNPcmlOKOyp4OkeTYXONEYzpesoWaM5Gv0HtceYF4u9vXTOTeUBZoVQWloww8TDw/Zcuw4
0dY8BQAbHcHszgjD53XhNWMjnK6tZn6oBRrnXxAO1fZDsTe+hJHGdzEEWZe8F2DG27x2TCfDHtli
YfkTfrDIRUkf+7hKjJNIzxfNHaUPs7kJq1WtkAbi1AAwrxyulsH5gT9EmGXMEtkzu09v9zKSYMwd
7xCZxT0M7sXr5eTp3VDOmCqBHHCqujbtDOuZDQD9bPAClj2k8BiEq7XLljFEttMecoHQ8Yp3izOS
P+WrNdUQM7EFvUhXWjlffFruNmoJdsDhKqlo6KospiMITf/Oo6HxzzlKWJArre5MGt7/KCze2Kcx
08EL5YZQBpV/FiLIpt5PxigfODroMOH92TYQ7s6/ra+c/uZbAPtKUoBOmFvVSFZqWmZPfFioGkP/
eP5dFcPCvSJ6q7a/XSReggrcNatr4SDXRyjJDhgoA2Bf0pdr2cIo+9Shj08nMHj6OzSmHM226tjn
JZ3BDRtvFHV73i4R9wrM8RX+A97EnWh5PuUgbEZ2rUhgrVOBPpXODd/nFI1l3jz3KsF/jqZZpmI5
HTpCbuctXcASsDz0XJrVGcWUo5nFv93erXR2COcQ4hwx0I90ocFD7OzZRg8ofEwOpolv5XvrQ6x6
EGAFLEeHSPEFt48F8SdygIktLm1vOe1SPoYPsz3vRXIMtizgq0z18Wpma6uoZrLiwxXalfGoYrKJ
ILZkKERKTyaH7Jc10JnN6wgiictmeAfuyl+qtb44XHiSGGLMS3x1Uc0FLWtBnMK6xB6ZR6eei5/E
w16mg62RZfDj5Kna57ynBqWHowCsrH450VOH6HiN2WqiNpKOBLgawsBFomTljr4YD0e2ai6uh3IG
YIHwXOJceNjeiBHct+hNjXTV8vm1lem9t1uTetK4GDAmT3y0Zb9hhx/oTN+vsTex+NCYszzwpKrP
zTXaMNZpJgWwc8gme5LqpPGJ1R3L5HJQEndkRGckL0lljb8Y2j8H6iwvY+YNSs3xRFmPM+nbo4HC
rc9J4pMSA6ve5siQhexz/KlCyG2gHPOwH2N0KVjnxtq5gG7kXhMdGqUQ9YJvRVcLLmU1HsK7Wqxd
GwFlm5ZEB1XnwmcHju7QK+4Fjy3FxaW8hOytv3WfhwnVmn3FPoh7bYjsj9IqKWDMD3yxipw1to9H
40zjogGKGxdxkJttqiCFWYMu7J03+rhM+X+2GllYtlUK/bg4kmSix6hlnXwvOIZvz01QdIiq3eBp
zmrex2/zTsFhUI0ZbaEsZKIGZRn+O0tF79Z8MKWZ0SvacoCIRr8Uhuv6va7MOhOoSMQzkAU27uCf
zO1XfDNXosAULRca+Xb2iaW/WjxPIK8WeOy+Bvmb2+29T/GgJCenNbRPoA3PmRWaqw4GsIbHbGtg
hRs9C76y2la+YtU02AQcvGWRQ+li3Y9oqVTFmn91/i0zrCvINf6QyuZHuadK71nDoilXXrWROCVp
5IHn6QuYjcFIdSbzYVWhRk8P/kBlWEb7CSiBi0D7OqwJN5QLdUOe10g5qdmiWRWGbfFDY1nFumxa
fSHqojJSDXEamsRlSIci5Ofsy1c8YmOcybHUYwaajYhaL9pkdnWwlm1klPHEW7qRJD++C0J5p0vO
7JyFSb63xWTqaRILF7atBwn7BRQLxoKlf7BlxTwhCfoKcthPAjcYkIho6YXJ5zGMeeJPmVg3DWXB
n4omEmThBtkOInVShCj1wPgT9GpAR/9lgrLq97dIwdDQ8d0vgmy3eNP0QMVoZAaywWj7+lczAgL0
+S9RHqzZtVuHlgqGz2mWcj3SAaS5qK4P3BaQEOHxd6+CiwUWOGvh2SGfDPIIikNerce5Wl9hWzIb
XHlBdlVPxhoah6VfQhL3U5qDNATy1c2CM/SfNu2KTj1joAQkhY5/yiCiNKmJfLynTIRffuSM2OVa
yZGLlYdJQd/gOc3wSM8tvVVmGzg/uOU/5y0NcoqVhhVLE86cVIvhvN7ek8iyK9bRbFO1TMRly5Sk
jbV4Cq8gb+0r9pezU1mjvaHay6eqLZ4aEwQ4zaeON4viJASzC6IV6MxcInP6iA+4XlkPo3gXWR32
mPXrVqFRtUWV5V2rGlA7u/TWNXVyrigyfOcS2JyxacJf+MUM/EdudXakun7lzMNM4KHqo3VhbEIl
2l15J5cxhuh5gzD7s2c6iARUUmJqTekZtjW581MwqiC4FGBWeGIWBNCBiy3ezGkzalKvb8qYJYUb
PXSVaAwNKsnApE9yy/fy87PDAx6PCLJKQgeyMY35wpWqhM0hFoMeK83+lRDgnih/36CKtsS0UmZu
TERQAy4ouJQ0H3OeYbUao8MGBjUW51m1U2elcevUVtLMoMNPQlGHkrgH2lQvNgqrcOgn+jxK1mdL
eH+pe3X56aZU+pcDLZJii3iyII3xz9qgGCY7UVXxes9C1mvB5KRrZY+i2dNliChTur+KM0zuZjbD
eZD793R8mWy77vSuHgR5MHngaRqPRh3TchaB3d0fmGCyp86dicLYUBBM8J3tZ2kTZmvC+b7UC8ll
IvZVgpf8PAZAQWb7Fa0366vNgoE2BJqB9F1ctXHhYjdy+MjGwyf/bqQbbLIHwUfg9ysidmoXRK+E
2xKdQ793+YcVJmoQHzAX6sTPs/ZSJmA457j+ccyLbvQJ77c+hq4YE2xPIgVpOn/SSHfX8NzxAjMI
mtMBIaF1umZJwwPRrkiMSuIQHUgZ4Mk3POMEO3Zq1NgtY/Jay/jWBgbIDcFZXyYMzFAWkmj0U7b5
hxoH+y7SNqVtqhcTQhlCng4RDGc7BWNmNrEUoHhlSuPN2w1y9Eyns94fvSLBJ7LolrxlDXn1iQQ/
dMlu+RFu6fB5L9K/iYGAE4BKkr/bhyyA5tKji3u7Hj5yLRSdfNNMvfh7IfC4hGCMS8/eN/UlscHf
KpV+Bc/ntkfU49csqjhgeIQy89bRvMcw6h9pbaDlm6ilbwsbx7aMbTcdnF0K9dMnO1Rdrb8X1i6V
6t1kbweS1EB+/Gxyn60pUeMTwNaQXWLyqWe1qRzLF/Q0V+qHjd/RngVPi8yg7XXmcDNuuf/zw184
OQsOnz4t65CFrQNKdl2qy41S5nJw7z2DjyjPZUdFnm081cI2iiVCObhNPf7lHY7xe7w+mJYXceCt
UrxwUQ6IPO1ZQqvYr+cwfXmM+li4gGmFB2EtxL2tG0f2i4IOduhYWCdiO8TxJmmCzLlqr83xn0JZ
AZ0V6ZRrD+8b282r7Bh9gbE07ZCL/UGXIHt7t47eCXMlaqGLeXSsBOVLJ9rQqeiSnj6sXGoV9OzD
JpnlWjqmcOhLp6tIaWjRoYbfBiPGU6qNzrc88dcleg6a1srgzNnF2tqjOs8RA64hUgs8hl78r7o3
i8ZIKhOZ6IJyQGHX3rHo+2LImXYvVa7ELbapnZs+muz7ePUg+Rt4CP2HeUMLSujhHjbPtYWbPt7D
wt2e+e4cP6oQgmUFTQLTuZ9t7GHHtKgIwQBkz0L48r2u0Ckvd+YOpfQovDuFdSJDufBuBGtP9hLI
jJwfZ3qz0N5jalUsExFd8wFCFGPJU4i6tfUnYy6D2KZ7YR/F6VESx2vk2kwRzWIJc9UcFpwH148Y
LMOSZemLb5QekEqQvVsvCV+YgVZNMvPgpwAvn5s9Xc6FkMTFqmt5c9JR3Dyv63bRegjMurkz2rzb
oOJIWizSCaTMe2dxVqg9+W9isWa/Z0F54qfgD5TcWvxG7UKPO2BmJVBoQ+H/zx68nb8hB78LhajN
Gtc7OW8y67iZKvGpBk9Lf0K0BpNpKoGXNFcFbKup/PR6UR0H115KyqRr8ed8rUJRnVdgPejgAuFU
wxx07bZdjKMn5owY/6t1AlyXYDIyDImwZPMxMy1qzRjW9UWH2+2QQGlcgQkZV0vW0wGx1rXXYe2i
6wRkags4RwLNcSdBXk2C5eplHC22AlEDU3WXWKwzfEk6Y+gis1WLNvMkSoa87fiZ2SI5rtrI1ZuC
KsdheSg//xlRl61A5/MSLPCUFDLMmhtApNvJuwI+0JJSHx19K/rtP1a3tV5zeERhDnr/QLcPe/iT
XArgvF8FWakfG++EwskoDB9j0LiqkO1peM5SqCbSF8XDhCM59rGfEFn47UOO5/wQvOHfOo7bCFlx
QyGNkgZRuiN04XqcpTkSYrdIQMz0MGHKidREfyAOaOys4yV09+t0lxaYf7zVrgr4LUW+IrPtVSIb
2kGhyTlNugkkMGKnvTHJE3f2lUflhtzB9Rj3bDqLPhzfP/FsSe8R/36ZnGcAj5zsU42qHRxOrfs2
mllXq3qeeX9YLOqzvN6M4CgTUiOjtqvPtQonckQPqlj/mionOToPNRgEsiNE53TwNWC1h7J3buIr
evOfRMKMla0WbCAZES4c5afEHN0g1LCDG9bCn1WWqrFz22sb0Tym+OsrIEb4cRhazFnj+AY5oBMZ
J8SOKmojeGKS4JHdLBEsAFMxgRiNH1+GVlWfTG22pNlSpdYk7sx/PTr/FrpqrqKHdyi1qNjghy3o
W4pQG3GBZgOVRt2uUQHyhjxMwYuDnMGiSoXAGMMsH4RGOtZS3dAiIu1aVnyl5R52X4r1WUzaaNnh
w3Qdqlmzx1/3K/rLn2NyKLqbPeCyhMSuDU5BBHyBUdxzyyyshAWUPZWjGk6Q7WiFptSL2jjeTPUT
icHNhIEmNkgPLGjJS7UPLnWmto58vqfwHF7lcFZ5RL8RDPTKpDnHPZ8FX2r5GP8P3ENOsPCk08Y1
tWtkOWIGUaKAnxMLEV5FhAnfOytgU/z0ZSCVI16KeR/7hhxmtX2Z7uLz8SSucRDmAbRLpyMhAWTA
8TxCskZCO7JBGLOv39SaR6xRDqRRUXOQrvtZhAkxsfo3B4rciI60JD0SbN0wqVyv3IiPajadGy0o
DyOCWf8uCx8BhKDTR0jRttrn8UsLTgOy0s063KvKEUAnd34usgvWxolpNqsatVwjsgTV8kZag092
u+TTv5PFZCreGk1NYuts0bd7YuVZ1pNPe9OLdQXCh31cLZzivQJRH2T0pMPXQKF9uicHXdcPd4nZ
p6lkcDFOpTawn6m1wUXH9++HdZAO/6eEf1HOL47pUdPuaqkAyO0slIePwZDohsCVBUB7UTqs3nKr
jyn2X+tWB8UtceHNn87T7VNDoV35mXFWJasdnYaeqEi4ueDoRMrBhQVuOkBFQFjjGXxEFaFKGxiY
HJsxKYYaj09AMI3zk0xHEbDpTv4wPRLamJZnhVG9wx1t6SbL8vv9MecvPNM56tTUO5+/QknXLHB5
6oX+9+rza+PEgCOm8q0kgndkmLSdshh4y0RGC0qoWw+FzcSsS/SgQICaCJA/p8tmAxxfN5l9/VDj
gvFSmjHHRpxsELjiJaYe9WcHUx8Af8A/PJFD2Q4Z7N/s3rnXXtfluaMBodRxymTJdBgASRW6f8r3
qjy6AFNxCxNWyEuQncqqy64gGeJyyn9fiVXM0YYMXUB8sGsx6JsH8KTBxQDeJ9lYUnwMbFCXDJPZ
O49j4FCIUOAe93IsIGccUXNwPglRrAc8WTHp9SDmGlq2Sf8zOuUjlQ48Nao4FXfhDc63d3Gk+Uj5
yMhdE2/ZdyGG1JxiBTbaFjBNPSNbvFr1L4AWQnWK1heDNEiMYX40e7SI+ulMoAzDlmmYLj9pn6eV
ygpwv9c2y1T1/2DueYde5BP+aprKepZJ9qz1Eg4jAuRGPO65I9xmlhu8641IvdmjshAO4coStCD4
NWkaUoPLCT8RgSvGGRtYYs5A79ZBCkC04H4gmQNyQ3Zw2riLb/Q6mr4zIW9Mi4RS68zcNz1G90wH
TbZV7vHdywKKxCSqqmrhRYpo7Ifp4aQVCS7aIcQAU2GGrsKn+hHFKADD/P7tSUUmvsoZaxTi46cy
y/sn1V8/xadT/Dgw3LXL3bVpGCM4SK9fqVSgwUxmCvmH277EMCjaR/rD2Sj7KXcEkznHwVAAbtOA
I4idsUxqJ4JcTpSPMV25mIwdRoZQ05s64YH6n6DwFeB7UbK9/EnsfA8/cS3jJOBkozLGRlit5Hp4
ESlVQx4QgaFZ4gdE8H8u3v60wjrqb7N3Ht8y8iX8+eq0iBEyu9T/qwQtwr6v/aU4hZycUzsZt9uJ
r1jJL6u+yIR3IZ9ks09E7KY62RxbJtKuGza7q981vhxh66nGr2q8lfwqtAwn5dvdHiHoZwY1RcHA
Dx7PoucHZs+3SMkbFb6vBH1AvvlFKk+AXL0HYi0lL47lGAe0FJc79IYdn98JI/yl1gmYkuCTnWeL
6oDYfT9LuHZrAy9R5QVibeZQ7ktUPxjd8O3zPAdsIPKPX/W2we7Dl693MBifD21DKOLWb2Wc0RFj
ObWBV94pa/9eX8k3wuelmuUz84JqRBjChiywO7dmHiXyXYxCQ6Gip3qCG+qT5k0WH3LbLIPw8rm2
4H9Q3ry+5K/SPsAvzvODL+ybm0jSE3Vb4eNWEOr/9q0y4LEiOlfgL04tOKEhm0AoLgLYOZowjpcX
mTIR0IcJd5TuBDwaViSwxFPIZHvckPEPSN/Jl/K9z4/VlrRkqScsaMhRJLDSvCpwkZ1PYY+Fv1dm
6trkly70N6sH0aEYM46mRbkX18HGmWrwvzu3vFsxwh3cT8KX9/rNTm65ut+sMWLj52ec29lIes+v
tWRSI5yXvTWluFLW5nLDsLYTIfqbu56y17NPaBggZFplaTnziXm9OkJWCy5XiGuDfSSEBWbz/YV5
HgkErFdvoVB2GNjKghDPnB1O6X5Ji8RYPAMJzjT/zfDrumxTFUpVtR6ZFbdFUET38QNDY6MxX7R7
fuHAK0haB8TRhbvxOsfMd+uqfNK6lJyhzdxxfGRNZZmS/zULp6RkL+7wC/222iGnAB0eTRRowP+g
2F9uF1s7XdGRUO7BZ+iCBs/lOJNMs3QrdUPShDTjLZawgK07N4nCQuuKLpZzRDHc/mBFRuW+yjSe
tqIAy+muuCgZiIN/ZOeP5AIS0fXEmEC4EEisjl2Hcur1d5HbROeiqyqJSs/47nyw95wv3Lonszm+
DoNs6Cr4hr5LFBym2i9c5DFqLutmzvpvpFulm+61CsjRZQ6dSgYFtUaqAggrTML/bQxx9gcmDmhZ
sFG6uYFn7CcvLyx2R4OitqPeMfLFqYsk61jIfWr4oI+zNo5QTJkrE+Qj22Ld2JNqfuIuXEfNXH8I
wX9YxUKXdF8nugzOsZoZeG4acqTLaGPGKJ9GwSc1PxaW6x+Y6WV9OfGhBj8pdDdeuIilANwIOtzy
AMBv6LmIOV3IsHemX+/+LRRDbHt7hqmIPimcXinJu7Cj5MPhf5zwlOSoPXygkktzwCJCbIEsUmYu
nB+/dJ+OwMX8Kl9R7Qnzns/8j+mpGVcJd1IIRtqUruG9WHPiAncX0QtoPCAfqEzwJAyOYqXW9gGC
885eBQnZY+p+VhXUuH8zhGT0Jl/6T7npowH6EzR2UUXsj+n1zEo3ZnUbgMc0s6CVWU62V72DPr6b
+rxhGt+Q8sgdYHVVIN0eA5SMMFNrc8iotNPMcU6FLmiwcF/gQRy+E2tqcWQGvcjy7e2y3N4uVB4a
CkmgR9onoP6GG1P2mwkbjQITe+MJpHWCI3PsAqoNAdDyFVQfo3QEtvjKV00mfscHJ+GmzQX4QKTX
fsTUChFJoh2BntWBqrGVuGuwsvfeX73rDeQ3I0Kc/CSM25fLaTrmWCeJZwKrqoK1ZAzbEQydfLHW
1Ju4FosgXXnJsV4LTtDSp6w3c1O9tR5JoNu1+ZrepaX86wlT5t4b7/RiN9NR17L3v7ejLa692Y7X
W6iYlG5WUkkLDfE5kOcH8Mm77cIqu2r4OKYUOA2hf2TZ/zwpWFi2ujXmVfeYVlXYTgFUaiNmMFU8
T4lGnE9Bp7I6XfCO059pRrPi7XYEbfpnohuzeh7NEdXEy8/FcDJwHSqzUdupZPWrFY5o5lv7tY8k
FacRSNvdRHyJ5O8EwAVqs46i/cO3Xqkhd6IZR//ZEz5dSCMiR6WojEyaNSCy42dNVtJqhwybroyr
e0zqRFfUc0ledUZG2i0MKNPIhsDPD2yQ2ZYVrtOd0B16ZtK/3fXnjhh6pna7y2Q8G7AmFzT9Hsch
EhS04nGjKHbUigIzBfwDWTCHVBZEtON6tkrTkyYo/RgZ9newp4QK2B4dn6OdgoOVHUmGcMTPVpVR
E1JY+TBCijDmWDCKPPvjfbfhBryZQvsLQacuTyh7b3YblAJ0Ca4673kY4HXOHT9TioZm6ZBjX15i
LvJ/XE1T2Ia5KQneFGGVTO5wAkMaEr3YpwzDkeCboUkv9ERrLpJdN8Hf6POxSMx4EJXdW39ms7TI
ay/UTlDqma7esV+YlPNOX/oi9D+ACzeuFvaBN02gGM3EGAgsBzHigCy5ZV7x9ENO+d+ZY4psMCpY
87Zpq0yot18GIyDCrCBLqSvl+Wc2KhhQi42H1PebezlmtnETeFf2PLAMp2xzjAlnCA5HNE1LGnm2
r/DVgI4rt50Y5ukt087p0lU1g8dtaui137UKjGkghA0EFQECg+Bu/MmcmpEEtp6cW+8q1bJWaIVk
fsfeE14+1dAuA/LR6lKwbjeQzbmQDbr9C4cE30mNqpU9bmjas5JS/LvK6pFLMFhrAcLP1Rq+4ZN4
W7nlCUtJOouZLzyIvDGYV4Ov0jjzf16aAnrZpwwbLdOUVyc70ZTphgTm27eF2etiZ9pJmSSwvTaL
DYCk0ffAQWc81niGW1xzegvHDu1UGRNwnuB0yyEZeANO/GsW//yC9HsNfWHunezY1XrEANRKFCmP
oYB8KG7XAHwCIekNHJEW7qupHwIQmOrcXz4RKwhifnzJUfct8O8SkRF8QT3recsBdWAI713RQXvF
2If1+IY/ivbM47tWi++Km5ywmoBT049bLKhoAZh8Q5idCvD1hutSkRrRfmbAI8w8sss5A3VBxv8U
TKYzXvTfeHMR9UjhbythaSpmG7uqOTMVSoneHLun/op0xElhwhOx6GM3oNxGj+mm49EBBWnX/aGd
AbByqZl6u1JxPth7QkcEuu6hAILpAMrNJ7XJqCb/RqkVhrdTadwadP6A6JhwnKxqQuFsG0OfMAdI
COyyocktC0n6m77wE9fAjThsADsupVWFRRpxI1wVMFGc09s/CrZOIfHh9hlAgaUI2kNBL3rUYXox
LjyvFKvlgqxHI/KT+rzPzTrqvSMgimCygcpmKBPv8laIw1bw2cCr6xon1LVEwVRskEaPUYQxm1g6
dORpd+ag7i61eM4TDvdW1khvIXU3YSuyhbxhq/Nx3cIN2jIfH8dQ/Ht/7OW5u1F7vRK4s73t/tjJ
kJA3D6+vTUUz50A9ko9AaSZCLcCOQNh+LFvR4CV++Nn+/XXMjrsYP8SUoPIH/fIL43cKBOq3tWjK
1OhfRtY8qT5+OI1VFadVIP4D3MKuc7Y20gCXeANJe24HXgCVAnB5+eHksDMFwvMLbNE1a0Z5YNeQ
5HuFmUdtPaztHdjmEeL1AFUea6P6BkoRpeprUvSrwzCgpZ2ZETiZJlon6T6Tbi6n53UfVGV33py2
HBXtRyjfmBhNgZ03I51SOURALuevW/gaKBiAP6iOkBLG1YUUZdAyNzbjh31Qgpy0fQzmjni0XNU/
6jQBvhDKtmAiP+81HXbE/ZJoIr03PQvOdTa5Nv15gaXlzE5Rfb5CUQAZd6WUqcFiM4lkdVKCwtq/
K99XXY3FiY6PH/4HZKWUe5xButr5VteMSpqXSwa5ps1iaDV4+CQIFq71THpeqlPFoYmXFMv7aw+e
FYHOY9w8Qe3MzgVZVsehLr9CPVd5yow+nBK6iFFGy566OUbmyfmVwFsSEV5V/1wTjKQRBfCLLoa8
ih+4RFMpRpqLGw+p/UKucASXyOGv5KZZang9iQo7kbaJ/mVXPiDAdEku6i1EB0xte8HKfWeLp7G2
NAG0rfAsrEGkQyh1idV6hFl/etR37Gs5zHK/UepbcjlbGHlyHFo9IxRJgk8rLOkxVl3+N9OHA+c4
BsD7Ow9wfRJQoTn8rW0HHWs4D+j6Z4sDncMveq9FKLb0c4MDh0BGPsA0XmjHYI5/1+JzbXuQtHW8
44TGnqeX3VDO9oDgBvj4lgNI2C/DgqGgtjGWnhxVtumsFeUZuuu/CC9GsbRJNJ1QMxxe+Z2jXGs0
hX6iz62rxnFogquuj/xGH2Gosh0sAf+/KegagWHkfqL0Bg+eePpAC2NGPzqMBJLRNT3T0tIyECGJ
7moI+zBPVngZdK98Zh5hIACD4lsPFshRAIoxFOQAEF7i7Px9NLq/9snYeiH3HhWd9gnQcohkJAWs
tg82jvDEmGvgnCjtPdBNGkOaCIvKxaGvkOWnWhqD9SGg4Rx334qQN5P4von5yANQdTzg0ilQe43T
qWCSrAV69i4+N+oCDwDOSD1xAWO00jzaVzGfyDhhC/0cCYvkYPZCuz3xrsYiRK74Rr7OX1qW7R9S
CJr3BySxpJzakDizZnUtyhaDJzP6jMkFcf1u1X8KCyr8ctrcgmNX5PwfEli18Pn786lHPRgeJv7H
fFQi6aBbgdtNETQpQKfHFmM6CHeduDRf18Cl2GDlFD+XZZmpFk5jQHO0hnynh9e2bG6G5jiSPMwL
ZinGKPaGrNU1A5FQUteijybnVGBuzHypis1EuJ4HHfuc4HK55cQLPRMp445gNirBVvPEMtlztuHn
fvCFKS9AeR5GmCkcicbsqZ92NVzDpZdR1Q9dfcUzG/zkKOFDC3c34XqQhWqF+3kJxZgd6F3bQAI6
hG4/cXh7Tqq8oufEQZd++tupVUaAX+KUhvEedMqGFEKVgeax67HY4wRcCh0Xevwy5ZDGigJ+4VYo
puFTB1IfPH02kYt9AOx1IHsuN1JEN/nwOEXyD24XPb2bKoF0StzpHuz4GeZWajJVB33UUihFS56c
lzfwq+Ywn/gBcgZQNlDxp/dT2W2BvcjfvRDEcOHpzEQoEGpMQm5SPJkBQcF88o8HNgkk7dhR33+O
xA4sHwYpizRl1iylf2P6483KonkRYRW0B3JDi/sp5Z/jtERqQf91b915/jvxQdi03GfZ6PoEmIT3
1NCgcN4vbsS/2V2WMOHpEgxt1drmp66Ljx3byWC1KFtVFzwy8fgmc+82iPb2LR+VA4NRV7BZm78S
ltqlQCTKl6Ths+iPr1wrbiO6sjb+5pBxw2SJD/WOtuboqiaMzhKZxcm6o9faPq+itimKc5u9llqM
KiEeUEko325GErA1k5DXm6sqoLPy0e5l7kqbYUjRJEX35H0ku70zsBq7xDlBeHG5JlONhAzVfxE7
V45SK1CzVMVpL+/kMiEKtvimAu2yGtQBtdCrs7rvHmGHSF67ZB7a9E4R+yJ6SwDTFwvitQLe1VdR
z45MGY8aTt393lzkJU8Z9MzIOrxY1SfICQ5jP/7ABf/byJ9SyC8hKNl3ei+Ut+Bj3bg7FuXq6jzM
QjcqmugBV9Lb6ycKloMDtusiLvQZBhzh6TPs5uw4wW1VKEaiWwm6PuJA6hwUS6d6dmZ5yrSC7Wfc
js3m2ISwRUj1J57gkSG3FvuFIGXtvuROsnqggXGVwJv0DEcu7yjh7W9IMH7+PwI2U42K1O0+Dxci
S+j2Gn6EowHr6MpkrU2X0+Oykv4StZ0yJI1gMD9YCb0c/BXZUPAf/Uu1UnFrcDH+SKVymZev0ybd
wlALuKzP1TWsQIic3TFdJaFozB+Ko6uaEFGbY5w0Dyd9kHfkJROCT7np7jP0AjMPjvIQkQsb2rat
JHv9yBuXK90lN950m1bFBRQCuadP4Iwq37qyl3iklMGhiFWS9MEtfbjBT0fzjs7avic7XI0ixWe9
qkGFmKoJeBm6h+r38LBALUsSWvtepPH4zaX8RBPnX2+d/ZBL44Ahdq2E50X+ES1SqqpEYGBisGHR
rG4Kc/VCoRRbvN9OCdxKhDD7GuYTcrfqi5NrxW8mosR6yQH6E828KaM84MYcLIGN1pZb81+1ism7
waH1JcQMkX1wXXOMORRV0lA8Rww2p/V4K+Fc3mWb7rnorQ0PYJvW7xdfHkDP5sXuZ9dgPZexeENy
5mj99R6xh/oY12hBD9NyskxTXfzFTW2dYwKDS7lqVhkRgVqOhnxC96jLJWGJavfj0xSsibdnrjt6
w7lBS/chov0pILUW/BREY/q3yC9Cg4hi1DYueTp1Gacr8cTkTewZtXXO+Vs3QZJbRZAkF3/CjSIm
9aqHvE9TRuCRuV63IFCyJfOgh7y9X1/WyPB/h4FoE2316qd7VhgeYkt/0S+uCXIP6GgoJAtiDUK6
y2/7CDPGXF7rK7m7hWK5gk5l/idWvLDJFa8SRuyElqjpcTXRG/uanMATNUoQTr/qqaNADvJotmyl
7gocI4Kkxq7kZwphD2LM1ixzPZP4+iHSiXTOuFzcG8HIbUBaz8KweEKKxeGaJatlX+GiBjhQLpHy
htt8nB8kunUD5TkoXilyULz6I7sohD+RnKJKLHen4bpqm4S2mYc/f4PvYnmDC5DpYUbmr5QfQ7TT
3jISGB2vRGvktC2oQZz5pHxZB4XUzP7SEe6voz0pddd+wtmCQuefJd/nvxqKlfW7l2uBJK2E3uWp
ySE41Rsb9ZLmUY3x/N1gwaKpqS9FOR1y/i28Q/7VQdXAi2erZksAnLBV8sakmwZbZbDszlT37XMg
DFVIRqRVu3Kl8g8LmHckfaaUB1aTe3AArFjzJE04K/xrOZROg1teLlQfBjisAQzSgYcPuISl52Yu
wPmyB1KTaP1pCN6Ee0Jy8glUu03BUR2LIxfGS2p9z5I2aMPu7yWlWYbbsBH/5S8YpD9B7b3MTaWh
ljjGzJG3JbEE4yTWCZWuQ8y8dBfRl+NmzhTqnFoFE3am2csUtkD+Czzbf6ZANmu7+/RDiCrue96N
h4cAjlnyunACxwGrq7i9T1Qhly2K8NJTjyhCajlpFtFfJMn0D7mjh78hj74UH8UG6GRK1bJAbv77
8ZCTekG7PiDj4VbD87pRfBSVlrywzc2zdZlQ50qBdKaEOwsR0WJ3FaOKxbQ941xXQQ1Q76uTh4SC
rTarCwpeIONm6V28V49ipgtnCyNi3Gh3MgG9cIew3m6W4/9w5QUsLPStWodBFvK4dNxSGdFUIUZi
rqrq8awxG6BA4elaipW9VtHYoqyksPezaNNGNRLIr3hImfMB0bGYwS8BN4ecyTKJnMoTeSYXB2e7
8GzLKVT+5IRO935PfSs9rIg8G+9jG6kOPujoZWNeun3XTAqKHPMvdXt7BtZ6V7vnrKU75oPYh7mc
pUoTMF8EJfg7hgbeqH8Pn3wXUU3z7ow1O+KvTu8bPjehBTp7/HZxjMIHEayVCPe97jg4dcvM3N0Q
gfkrCuz3W721M72sK8L6FzpaGq+HwlFasdo0BTtZjwLheEFYrhFU26Zzpz0NoLUUI/EcWwb6oVY7
NLgrJ+DzVDffrQ6mXWWeq/57dFzeXcE2Y+0n+bkZSwRzC391Nu4xjdssQGpjmC1ndgLme8hYw8mO
CHLkVanC7IGQIfg5z7o+FB/efYtXco1+NjMupfmNoBE2AGXOl7eoDMVNi6uQ7QvUbqYxMuM2qkJ3
nZUUjQNJOdyEWVWwQ6VSuqeWHt4YKBYtJ+bspS3ZDVts6wWj30Lk8asp0I/0g9jJfKicYp6SvrBT
vlzbqdCQG8qhrlUt73vmWXPv2KPpx5+gH7ZUsFHRIYoaeNUxcSdiwPkfU1gi/5fDfnvcDb2t5u17
PvCogIqohE3fmHCUsRyYz75ivmNmWJe/LNr4jKvO7/UyDyeZ/bfucfd9BmZkip7RRR5EXdrVmLwG
VgtYhBTD4nAXzYMkFG1MNj5KELLgJxji8OzQDQ8LKkE5zJpcIwzan8osAkGLFBrAGGZsGQGPVsUl
qtjFph0FLDrsCotQMOA25E+7KMjnhdZoqS7oR1y01I+e+dNSF5GOtnf7mJja136c8GwwD1z2kr6a
Jgm8Azfj1zR09PxTbTZoVYmZm+EKDWUfa864/CxI0OhskGfnATIz9tCPc2Zu09j1BbGQFnBwfZgo
mCcXUS1cf2GPqIDhnJKsjOHyCUbO7B6FMc3XBsdPLD7WFyhAPTbTvbqFpqipbfzvj+rFAXnpT6js
/rkIacLnAt5+eRiEs3mg2TCbz/qcepzUVjGVh1lOw/9i2UwwWdp+1GV8P8UuhXxLbZGEKO9KyD8b
AieSKQKprmCxYTufY+ZqFiFjFZghF8RQPeb2a1FfiXv2sCqumlzXQvCO7ZhKfntr2xVe+aOJWTvU
3qteP5sKSpf11j+Q9dJ/NusKEegat68+QB092VKiuqhoVxnpBUw6JNPaEt80+Z3zYmO+/920i3xz
ORQkwl/bfBFoH5B2A2Tea0/7ZSTOXjvJsBa2+nCGlwaDDqFVZJ6Dvfg0J+E4IpzEHQII5jJOHqsY
xGJ22daCoURaEtB6MhTHZPPfaC5XDBi+XQpeOj55Exn4jF344d661PeGyCY2bJgKhISdtdRj8mV3
apIDwKINQD5c410azTi/PUXmFrAi943CUNCe7bT9NF9XwPdiYydd0J2I3aWY768gXwezQEQ+VuW0
Nsjd+cXQCw0F1rEjOaTv2w7UxS6PhtEiA43Vl9XvI+Y61d7KmXKIyylTkp5fsqaHWZx1tW5A/FWR
zGgdyQVb0sbuC75aeHnYUXLK34h4eLadDf4PRp4VlfUV/YDTKHPt3R4P429yo8ElAGVhdYXnwdip
wEKSeCYgNnqbZYz6DwSt1pK5bS7XeQz7HgldL4ahTsgqHKwdjSu9kh9aHGSCyT/LiYcmRkwe1hZf
A2ZcOrWVmHeZdLZbhgymJbDTZCjF3wCD5/iOghdvrfKDmJhPTbeTrpiBlZBPeVr57x4cd5nEsmDp
zHqjzkYSTAX1LYh3Lwqnj6Fe2ZbZPzwXRFM2ncxq0W8Jjmjr9wUsuLk8r+rwcrtORKIX0HuJGTJx
a9VC6aWPJxrnQzhZDnDygnAj4YpG52+YbkaeRYhOWtNRw9HwbbliuSUtD6bkNCK1ijca5cvMGowM
Loi2QT2PKJrNYEKXhwk9tmJJdktqtMCYJ5PV8xPC9g/57p1qfWbSqR3r0yEBrNa7JoG7s2QsBMIv
RrwP1HOIIvAnGghfyWEHoUZmeLhJCzY8Yav1pSJqqIzK1lR5aD3q4Sbtdg4B0Ub7juVZnmxi8Zok
l0O3Dsky+13NppHicnNbP1Y0EBh0+JH5/Bjr7wx1+JWpsJIpyslFLCdu9QREc6wHoXflWj5j/Mga
Tx1Y0uqlcC4Z/uBVC+xEUNiJtQ/rk0ojUUT0adUfaK9VIXUS5TmdPN4GM63pD1fNLEmbBbsXFFt2
+oyqGp6sYtK3HxrgvrvHM2984m6nv4S24TVbEfy0vvUDbqTY6Vnf+yKqDv9fvEHkkv6bnUboi0b6
N1jAcOJBDcUSafivdPWipaCKHy1GBJXm9kGZtdh/NNWiRKp4NWrXwgIkC3g2i4FHqgDWx/V6XPSX
uso4Aojxn5RAz5IGdtstXwJApcGd4gKhi9DUcWJ8/ZmPxI0QO8F5R4ObQs/D6pAoRil2Z7DJzeju
t1pFxpo1AbNipDYYwlESKHPtaR+lT2UTLSisyJ22RFumUh3yzzqne4WFWB6/pNSL+SOCijRT5yZ6
TE6IW0871aifRLYwv6AkTakJYrEoIRna7cDO2fGPahwnyney5PR6b1xYrtSmcS5uVB0kRDVWRsqn
DuBiqgGc1fP6LyniIz4ko2dukXxl3kqGYqxXmm7wQaAxP51DmxvmK6qHgZxprIbhuCdyNez2OPKO
8cjla8EL88aDxGPRKZqQQdYnTMHnESNerMB0xBFeHXjRwFsxoELOp2PQ9aqL+uY36pqph714o83Z
2fgTItStf2r9sSja1Ej0ylWnzd4U7FJaVZ8Q/6GU83bIvpLUn5Z0wxKioA9fkxuSHwD7QADz0C6K
myxufcydPUx3PDy816mN9RLk49xEbOiosh86ikPF5xAQ2C17RaaCq772TVWOiZV+MUC5AjKCYhuc
9MiULYIYyn5u1mmgDDF/UbTEhiWkIXYkVLxZePnHs0CvhJifZ82OpRqy7hFKj+maTEyet5WkVoqn
o8xcboNEH7z+uSAqHMuzTQzttc2UR0IIkQT6CEbdL2bxG3CcC6v9ATy+ydT34oqfHXC8FGQGOrOf
mOEgMHKtTSY6Fpi1gmdr9bS3C/BcdPRIQJwJSbV0zPnFWBCcKAtxttiypQWmapzMvEilu3HUabOW
NkfHpG8wIJJc4Yv2KnLWVfRMdf5LnUU8WtP1Rb15qEUfFXzdfCOGLeEEDV4kfrVsFq6i5eyIbznB
vvPW9fCxnFZv23aLTeZd4PNAz2Ims33InEvYLMNpq/MUOkuS3bOPSoO2/80GSTusqLIBsF5mjPuu
cxQqb+gFlwVBPJFP7lJx/xHi2usR3JE8wGtiEmWXZkHGEMotGKw43zE/CcPAZZruPGFUhh3/YiAT
G4XmCOxEGDmmpUjq4lHv9REBpPBnQ3Im7j0x53pMWKGQ8STaMMe6iFLxDEC1G1qneEi1/4U3EDo5
dmZamjROugdSS17ktd9XuKYRhT5ny/RD69I2b5grsyc0poVHaarmkZVb6hZSNJbNaqpstjC1H4fr
gpsRg6VUinbJLZ82/k03o3cXyao8EXYOAHQqf/4bUngHKly6ZOAuINl3mFrklLCVWrmEThP1Jarc
FqvGX5KOUzjfNHV5anj4MWnMhZHGJUfNe9hMhDtx8c+HjMqR/7O22PwOvlB2aG+gBMe8xLzF9la/
zlLywSxy/tqnQmDTSrD0IUzX5hr3WELnyIXOZlHtjHZBvjjXcTcHGe7zolKWFMBdSgi6YqKENk+i
f4U5Oq/tbEoreChqjzMbI9AhqEZeqfAaosjVRciGRSghG2kqq9AwknQQ0W1zUwThtp1W1gytpWd1
sADbBKOOq0PPl0zaJ0l5+TZ2eg3mz/4C0RavoUpKNn50MteETrJomtPOD56dYVZYihtBDugGfcN1
O3+G2x6bt3p70ad2oqTbZ8UJfWZ2oupMoTp9G/L+1E852fpFBTOA0PWaVD64bDV5QSb43uo2QjG6
rXR5KPa9xa6Ww1mlsCK2NinfU9LC40hMZwy6IFyYfYWT1fhHBE9fUbxd9waDC8+N75/tV4nMLHzG
TdCMD5QqFJuPrKrdVlc7NaZ+fQpdpTZL0X/OZUnt/WcPmp4CSjLQD6fcAUjwlLryBkb+j9hButww
yBeLVbj5RrlNjIJQ2IV1GNFed2Be9Ac9Sj8P9kcoC2LzSqP6+TG4WaZjVOd0HjhcHKs1Ri+TiGOy
nPyYhOhpamTGh4BWFU6THBM9qBpCXt0410ffIdGCBuiO0dNjb8wgwDIh7YKkIGZqERUbuwFGRXDh
vAbnHyC+x7TTQGYWzT1PGF9RgBchs6dRpKWg1GCAitMWkig4dYEkZSmT2r9/afeSvbB33itSZh/O
tdFzAdgzssdYueZe9d7uB7fshWLUiU1flEo3TzoEwSeL411c7KtRj2ghoLu5SpnMZXUsDRL1hIob
aBWUf992SKaUcYbDzbtyNShbQD0v6CGCqzHvZvj9K79QPsZK/5N1wFdMnmPB48z1Lbl0rPucpqmO
7mm82+JSr0xW4H4b5sWiACCtMTk0I0yp+olVQwJaIKgPHYRbIcPQvFi/LxBVdkdFK/+/c2qvoix8
ZDjux9IMc1kLlEhZsMdYvNEGTcAWZ9hqEDksFP7Qf0odtUDj+2Pl1mlPTbROBXVKd/RoaMlXdo5P
p9jozzmNdcC6bpCS1Tw5NzutdD+GCKBT56MS+La8R5EmYmG7UFyFFWOxTOAXiyD0QKQQ3/w+J8Bm
h3lhNp3xUsGTVvJCm5oNCA9/pn1MJnglgRgNbtwRKiNrEgAI5lZOGCJW/OxiFpIPdssJmu6R7pi2
Oc895R2V18+9qDWTN2VCY54DEzxGEfAuAKiK9F83fR+/UXJ64Wl/D/dj4OeD3p/9WzXFbMP05EFW
Hu7OI6mG6ONRLuH+J2uu4rs7R0O+Wezt0lcIefEYumjV57XoIHk2V9bf3xIbJUo1EhAQOEudD8gg
9ZhWft728cmAXWVw2bgNX6D098nzq/7aklh4FnFv8Wxo95AHi9alQit/JQ3vsSLg0XRF/Hyb14i/
a0KqFnrkUpvlbzVQRVBbPIznrEhwRhLazEuI3TeULNNozhE5e+SRfwmP+cKWEQpvnL8+X7RqkYG9
TZUvZkGI0gifeE8uHlV0bIOWo+Csn/KQ+dsg3qkjWT3NpWPekNnoH70/EXK+VA7OorKJ3C6+WrrC
HbfRkzuO/+wKDRIbVlsMrxDBFXNA3jKFvikjdjdTe/ntAiqotXkjSYp2amMOfjGQU6C/LxNSJFEf
IvSJVIhabSc/QIobObpHVI+k1mfPhBIeDl6Vsze4KUSxvIy9PKWdW8iH9HN7LNCV2Fbv1zBupWoN
r6CFDCdlIgnpbLQt09B2+G6nbKLKir7LMiat1+QNvdihxFWdsIDQr0l97t+B4VYLxRN7yDDk0mgo
r9ZFkgO9HeBOADwSuVeUnRWr+mno7mspv4VSaCPiALo5oZFcV3KZj1xnMAZdN18LSE/iP+pIAhCp
1iVizzaxByt21U4nHkxszzJ/PiUoY8tndsYexp2B1zUIz+M0NBMsfDnU+ga+r6FMPe16Rv9L9h97
bUnrAm7sST+AYQgFsrO4qyuypYh7bNnOOZWPgDxHMhd2LM2wCvGfKaDBemZTMtGH3h+e4NunLTBa
rnU7GjrwQ7X06arG671UIB45HAvnVbz4PaDFK9XYrHXUnefTgTeXceFNxuYaaR084GWgA5mGp2SU
9YKvGMLIAQnlDHT5NCg29vA5BSwSe1do19VT6BgPiEJZhTqngjhAc596kobgIKmUS2jx6ICYb7A4
tHgxc/VR6L6zyzBMGKN5b8WPCav2hkvBYMUbqR2CP2sgfm1zPx4eGCRuAOSa1FIiadSRP3VE8Ez7
0csLB8Zs6Q96RROEdw0ucKfkE4BZCWrMzmUJvoxPNauXF1MYQjBtHskvb7CQDNOykq+yxiNClGcY
ASvUnxZivSzD+mkXnG5vcqEnodDm+Ery5qJh+miRn8J2yZqjdN3UM5Op3r4Am67raLqMF85AEgtk
0iiYu+DYDQgEBStZUARN99wwTyUpmcENIhvzoHoAQInKw5g1gtMEh90MH5yjrF5UjQ9sE6GoSc/K
9+296OW45cWmC9Azhzdh0xgy4Wsyhb7HwqktWUT0nd/eml/w+bOyFa9oUwuvRC0J+sCaP+0jbZbv
6vvR94qmRwhMe83eviwi/EZ+0hkrlK2wlQjWBtqu9duo/ItNyIqqEDGgunIA+rLRwodv5k7r89pF
DHAQ8ZO+cHgMJppeylx4pj/JZT5LzO+siBDXT3L+sR9fL8vBkwewCwoSgu7neqKOIILV5XBHreH7
IguKA2erCpcRRT/+QBomm9uIUA9auIYUze80vmJvJPbRNxGeT0TRZRKkWSgpEv31cblm+zdYOI06
xvHb99uDQxfk/6qzjtZ+e9p00nmbVIVUbV56p2NS2SkOUiuEE3r1T/8J/gQFTHgS3OvxL6/T309s
4ROXYE5jdOcbKOX8DVcP7H+6C6nNqZC+KN9DARSBXR+kxuA08sCOS37v9FPycDRJWKjsWMoLP2Mh
2HPBeT7uMilLldRpKR/K/1f/g+nY3mhS6ztd9kcwl2c3Ff5x31RIhtO4Sk20+bNdt8+z1XL/32M+
3yhJgHKzJT5kAd3bwnqHr0SX1fSCwrys2yR5QYdtXipQxcuNOu+JuoGrwY+fS97Z3qlOog8wFdVC
3EE3cLFLdlQ75zU0xB4sYiKlIBDBbtxHaLw60k+BAIBgvR3pqwIUsxEN18fUppp/rTjIFLuF4Ezp
QdJJ8uvegsfYjXH+ZCdv8LoCBXRIqGg4F/77m8olEgi0WUlREJvSaV2oDBOsxwSz7KV16fdjkhqu
SHGzdnH7hecaRlpP1mL/3zOrv3EKjcdZbAChuZAU5KYYjCSh6VyK/vTg4I32Lx+NqjFRZA9W9eJF
qiw9z09G1oz2QLW91gGgt0TG0O2bfgayTP56RjGhmEV0Axz+ZaUcpnlOH35rg6xrhttijYYF9EZJ
vu/xTWkxUdt2b0cFEKswRvlpxyK1AZDZOzcz2MZ9WRG0shTCmPK7vPdjIPw2gYkZcdKK0avjuYsk
wu2sr7wEtTh+1GocGEBULxQcyvXlZy8RblOQsxWKT7/l7FyXFoIkCWB/DjgX7s7XGLaQYZMBO0f2
dxVzIeuvSq7Z+W7KtrUcXUyrzp3un1PFxa4nStnKz3qvAdn4ilQ495FgXzHXovtImPMf+L/Xjd32
Dsou6xhw3SXvU0QGMaWurqihgyz0ky2ML7Ukx4F7kCsDV4nka8pX88iGNaJv36jlVNvA6wn59bCw
7VFiAE765ZSSTXafMiE7ajCVdEGvf7uNNTW4zHng267PmOkr0mHAbb1ZenpjGJ90QFlVl4qS+KuT
jHXEJE67OYdYC+gnol2l8J8zIy+yPPlIqJjZAs2SNkDbUG7PRBMeeXDYNfMBn/alQx6gtGHht07z
wmEfM+HKTFrDnchA2nT7Jnz1DlhKMGpDCA1y1pTUT2zwTZQOJlpbQmQqHZRCxwEC9KqrCYBLZoaQ
nNXUTu1OOCVWn2WcdV18pGXLWX+ackSNa0jx3th84FYY0XVAqdmYU15tLa8MEcvL3oxFfCgKlJWf
1SX3fEfD1e/zySLyfCeQr4MVcfEbFd26CyRRBdnb++xTtQJaaa32NrEltCKamcDwBNKtsScXmtKB
KT33h4vB9DL8x2psQjJnKkqfiHBNqRlWj4erDO6tEomWMzlZrNiC+BBUuMYEAw/7r5i+pnpyYyiB
49YzFGX5XlH8uEeGX4a05hLv8x6WpJYYiumfsGyDw6R4V0hQsHpHMGIayEszwODBRKN6cBuFwho7
N2D3TvBaW6SvUvcKFMAvTsZYVt1dcAJGfp2taX9ArqnMz+4pihqwmhfVfhDfDoLE/Pf8Wkt88LuW
J66ZVrrJybxUuByMouOczbCdxWWtsbVMuzEdP18YItSi+y2U1zGazwjZd0A0PDlZQAvbRnwVaf0k
H6PeHBuozs6s568EanAqJMgzVIEGmTvUQ5WVYfnosej3UHKOxggV0h3+FnK7cxMzLwPPJ5t7sMFH
Pigm8B7Setl7QPe0Cp26gsokhLrgwu9sj6P0HFgwHTSfG8j22FRFfvrM6ICAkSRweT0S4br8ZNip
rk9vSx4fkGZpI+6jQgserQd4aUnmYejzX42VsSGq/6JJgi2PRmax9XSzad9QpPb62H4FFdDgmntB
WTRFT7+HVDyoxNrOR8zg0DUaBeJxtetAgy9KQM/oDcsOxEDD6sqcccxyw6Q9qtEN7H1CLttQXBso
qyZyUY79Xu7hWTnVhSokPkkwJ/rSEKzw/RK/JjYYMjyQW7lOzOsnwj+y/uS836kVKX1BuswgILOy
DRxxH/6Oyi4b7Pu6B4xwbqtG/U3QOYKNIgvk/KAZ+Sc5zK1u00j4LD+BwNeTYlr/Bm5abjsKpK4v
iQvv8yxymLZg/nSLZMB/+uy8W/DelxBlwhwG7l3EziMXrV1Rm5bw3O8E2f8cOpOqLM4oh+zW0Iej
bqHI8BvLzGA+Ttwp6wwCeudGbcivplDv1iUfSQPTnSgJ8TVQn/jE9eljbIN5qFeasl9NbczRgpLc
42sPsPxmbiFOBMGt+de/m3EEEW2Pf5D0qsxsC37vscXbzDFIj8hcsnc19cs4smXeaqN8ig3RSwpP
oZcBkBAHTv2L6/m1XrpUHs3jJTiFnZT1s1rQUp9eO3o1YGx8P+WRXz8GCPIkOVi7tb7adKihrNPk
7WJLbIT8fGQ7qiIHKKjL3a5IX3we7Sqa4/1Vy3rizmaUHRZqZuJnbm5xiH+SU0hlWYxM8YJnElZh
g8uV/n1AmT1huA64TeUJbg+4+51iZCyUiYcEJZ+qe7qsc6yJMzI0WUrtn/aDCVIunL1QyuG79iDz
BwDb3T4hT4dI7vQrPxHZfbGPX0yluRRL1XlircxAA+Ntz6AAl7IXBZA+0aN+rIzgSMcmZ7i+ym/s
cex/fJWzWWmspwop7D1QLHvJmVLgF19raJapfGW4oDuIgc04MPpIv/mQeTzmvHn3AcZx3DH6HeMm
XpSKPEoDV3Y5IlXGVP6lWoCjZBKgw6s/6+VgzSEvbCfG6fb2ygsLRG9jM1hboyGLxG3o2bUKjItS
JhA8jKio5QdWlHD2BjAB0BdHs0jxAYotwfCUjKL1T8eb/tN0EckhsnZimvR+rQQ0KQ6wGzVCPW4y
nENvs9VUDOdSAsoaBFwcDvKN+6QO7x38szVxrFXXffH8wyiLO7L2intgU695d62SN7Kx+/UrHjAd
z0tOXoYMp2CcHm6nl4hsD1ZMa/TEk6ZFRVbYFstshd3kR6Y3yS7bn2/XkswTiQMAjdzqHwBekA4S
pIfte8v4BuAtgvjdMt0/kl4eTqBK1UkNi3VrLhFyfu4FLLTOPB5pE/uq5LizuCYsS7XHf7Pfr2TG
xhvAvaD3ZgmSXB/83hIIq6LHyv8ZoHtQMopX2Q6U4qW1ioRGeCwlE/SntaQN86VUdNeSoMXM9x/h
gaL61qzPce+BE2SfABtRK3Y7r85ztVf1KZJokTBDhwyEtQpa7/N+U6lDDDxwAH1rm+2uzZkxGpk8
SrvIBdXCPa7M+4JByHioiLz92mi7dUvFt4xJjwxgTY3VuRq1QpnUYUTiarOJhyILro5nIAXlQ277
vLG2N7yF9LdFDYlE4uGPa7aT61TXC8+dq4urIXBsSts6sa3wfUOgwFNTfEpewHdbHvd2TvrO+Hnr
F4zbngNX7uQDbCkxBaiyL5/sAq2DB3KK0H/jNGhGymHq0TfzE5BKFrobXa2zfWoc0cdJfzX1tOG1
uZofkX3SM8sSYXzM0vGTY5cTI7DRmOr7kMAqrJfbRLmoaZdgTjsw7XRNrrAajHuLND6CConfi/xq
Aaq8x1zHuVOnh1d7g098oTAvfuMlkEWgfz/7Rr+27C8Adlc9sUsGdI8FtFf93hijPvTyD8ZllCEL
xmE5NtH2Yh2/bg2H+dXM4HFG4xPD2LSNhE9kmaqPbtp/4T5GUv3NK7+T7NxNrECpbMuFJnfyRQeW
V/ra2k3SbUn1Vlkfn6Nm9c3mt93R3ocJg8q2TdaSg6PMWA1iFYIboDc36XUuCVxCaoFA2O0wYxpk
bRnBC49f86ptLLCHMfWALXB1ew2PyYHJhIQ/E828h4W2WV0iqfiQ6FrH9H9ImRvU0eSv/vZMG/su
J1kh6FSFcmePtSdocrjAJb3OL+Cp2bJAqmsZYLSUnSxJJ9hqv6VJtVDb/dcvjLFCadBFRAdGlUQW
5hbtjdR3mvNpnlNcxTBKm5VsjygQOFgKKLpttzR3Wwnc9AfafcnCSNCVxwfu1RBM6ckwJlYc7lf+
BnHjdk85DUX4Md95jYJPa1i4VtjVCB2PsMCN2Or+v7dHS6cYU1Xbf/st1kFhI+/AuJZeQ40s2fZY
+hgXp2iV7RUpTKTi+COvVl4zoRE0tfYj3oe2fz23z/px9mhQyWkKQlhhpa0Pq8ukBrPFnfuXSWmO
nDR44dUpKws7G9PByGsvJoVCDmPBiLrrshjiCZ9pe30CHimDiTGgUNraAuj8FYFiaLqTGCFoOK0L
8g34TQxtK84fxc4fNyRvAbqyTcDFmCaGQqtNo+m/NPxeFWSnqAZ0orG1kfajjVAnGAEITfjv4LIU
Uyngp9e/r1rDTOJuWhACNd44Qo2ZbhuzQ71mhm/iqwIK9l6UqkA1PMCvDoTbjtX0YlULiH/nprwv
ynpISt80wz7I9DUFdQdjKQMvgD12PYfHH9pYPrrBIzYegUPYQ2T+4wzQmrmmy7O3D2SNkJBngTWu
w7cSUBgEQo7JOsTGxByyOKcq7TowmPrnzZnX6SvynnOED0RkGzd5ihVZsf8huMcIwciX15Pgnfh4
gEvsUOYIR1lKE/tEXSJFjbsoU6yOFVMF7m7+Y1F0IE7VlPFEw117+GyPoRH0KmSECwj8bSNyxNsT
9RKMD1DLR1zXTz1tljbUN0ntqpD/1Kj3RQ/qekHxIwW7BST17O4RCKRbAJlOxJDAqHR0hw+u1KCA
WeGBp2bsb2R3nW9IkGG4Lxtk2zO5fCaxYuzy2MiQYwa7Is0EWeSM4EKfiSDv0gHM7/xpt8RacDLa
DqaLSW3/K5NFpFGdAMITimxzBxLQPoWpi8XKgEKBfol1VFwpaIVc4R3IPWFefxAPLAyxoUaeh9T/
tylRdnkylV7FaUTfMMd/pKdS+px2GDrggXaseeEtVVnBDvgTZZE7RJTN38X2IxYz4E2Xc3hRugiy
Rp7DNcSRv/8ETLNVhs6mtWSJ13dkCVFqF+hvbjd3MHO7eZE8JBfilGJSZx75GvTaI6b3UZ+w8FC0
7eWNYttF3wyFdQ4qfrrPbRDI8VaAVGujjBP9/aB/j9F9Rv1eSKGfeKDtWnVt7ESu8nM6vEX+VCnv
OZIgELzlg3RD51Oo0xbYWUTuHhs+O70bYSn4TjPOWH/ORMrNDAjNV3FBAPRTgjJu1bMo1Ql5BeVj
UVBBJFSnWUMRCw0i1UsVRerntyBB0JzkuYEgWH3drwjdFuZxigs7Qa6+o6/TvUD0o99j+yEQYkm9
Y/2DYxyFtD2W56UPRTus89lXCSA9nYgN8zcFd+Wi7UO0q4PbhR8eEYjePOBqfRU55j0U7/lka/Hy
LcjRg2V3chUIIbT/wHEzztEnqWdpQRV8XHn/Yr20xK5NkiQPr5yCxNEJ75JQz3FnWI5s72xxEjJk
6c25Q8eEhYpN8tbOHKHkUO/f4y+VKBTuLfiBcDSkBFdhL/eCrKpddnsPgIeHyoQipB2xjwxps9R3
Md3jbLbAbcMA11ofqmfBNSYKvCRx9He/Z9Du0AdjaMmQF5IgGYxoInFMtAcFDdGRLOgz+lhUWPDl
U+J8YpK/tdJwEFGXNRr/w0tzGq4/DedcvdUHH+mSQKurZJbj7W6qFnPn91ebNuCpIHF78gyG5JP5
7qeSd10GUpMx/PaUoB+obWl5C/AIdOsQA0/JmQwkenHI2c6cQYcTo0nftuuAA9uyvXyPRmT1R0bh
0u3kT2CiFqnk0t//Nvp+ahFF5lCrrUf01MwSfrY3EDIj9KQMeABCkmH1TgCp2xhJwMlkolJGE7C/
YH32tXXiEE/EQWLpxEUUTKSp0R92OediPF5kar+/jTcmikOVHCHKb2ps6kSPKFQsOhzw+nG7Sxhk
Tj3SUcGuNtCC0yUd7L9ZDszoZOjF2fgWiZXFiQJTg6JHDOde13cafvdViH8A0QjPblnXfx8wiMzQ
Ft5YIsQTsiBjXuEIq6GmVC8eMGrD99ruQ2s4mUdQuBKAhg76DeEnfEVb5gOdJAg+loOEkHbnRISH
DXYpJXzH/LV8c+RqFMElWUgb9exxG8qBkC/TvB+YfYQVzCc4VP1eXURZbCOTPb1wWPDSpFRPCqia
/Xlley0bGsxKVKQVUyhmDpvDhrZ9j3uWhKHsR8qRFJ/PmlPaj94ukYliXmgbDKYIiFuabej3RKQu
gdT0557pL4CksFpO2oTXLWMxlnKqzbYBuqWxxRAh3vEtE4LaYbjtDz1/MLj9FbEqN/sufjbOTp8x
uah9eiq3HcQ6GuJYOZJvlRcRHN0cXG4293vQ3Bdz5AHip7A/aOyAgPqIur8WD58c5U9R5luV0it3
uBMxn1m56/eBjBmjjxktkP3go2JrdifPDkzm1iQiG+HWP3hUSB8Wp+Suy/JKY830XOd0EIXgQ0NV
INBmbmGs+K5XpMR5LnkWYitCFVxt+wWQMsktD1vtQCsix5fKnREWPD0EOdp3x62OmilWsj1FqGvV
gt55ukX3LFj8ArEL389BwOqP430bjkpB4urFE9Wlm0oX1hkTmJdjiBPyTl/k/PwisH24L6m87Px6
kxWS3YHt/1fDta8uNMFSoTxE3zhgCE8ldg00aRDiUWCdUW2RhgHhghJjA3JOmdKH85mTF+h/tIQ6
JomZ/zE9MbrjkCUAvABUhlkoo/4Vefj3hDcw8YtwMw2l9GOdKtaUEBAPen2atcI//hSfCFm4iFsj
IV7I+l5lZjn4VTp+jM7E4xmX6ZsQ6gtB57pcvATjbFsQpJFFSKfSSAEvD+uq5tnDIj9Hns3/OxB8
fq/hEQmk5NeiR2b9FEVmDfpaT8qPxjqWH6Sr7/KsscpTBadlbr4770KTWOZyk5Kp3DTLNKH1/lOe
l2dNzUVwsLPUhRfJBguiiWLgoFtyHw5VD02cTuJgzbj2/YSiVjZOGaDM69GQ0J2oCN/PrpgGwAEh
TPJDvgffELfDTGsJrEUT3g8Oq41B05AP3Nx9MVCn1IXZJF7isTvmwc0ufI+LAD+2iAUFvr/wFaXm
893pHaUS4SoqnGyELqX5gHn203BYz03Q5OqZLWwW2oi3xP/M6RgFcmvTKMku+wKVG03pK1jDppIs
WOlOCnypc2ebjgayEGobgaMx1je44GplzAa03BBj2FV0J6iRC1fkmVkpKHDBM5+b/vZqm12hFVlo
NB6V/l87eUWmk3ppINhjIC5Q4v+X9YWNAQFZTDy8SrQs3uohhiRbxI1nGvSHqOun/j+cXA+SDB2A
pVz1kiWw+iLu5CMZ18qZ9RtMTe2KZE0DwmV1R2d/DK3qLB+eNKHDd4hEe4Gebd/pKqJli5cFGjoI
PgFQrJQP5ZK/+4I0+IMliGnxMB9C+WwV4wnqesMHH8vmaS0rJ2K32HG4XKHatavbRnfvm4gEWL6y
ea+FckknRIUe0KNCgjRX/Xf3hf/+FsoT/eIeYkApqt5dzcn6rEgoXLDlMvhsv5xhvHTCf0Pf3Jk5
LL7WPUE2Pwye+QzLi8xc6v9pggKvOCgIBrYG5STXHfGnSiBcsLoPHMdoHg0KNsdMBYyN2BIH1V4V
rgaG+f4JXsnuwD6s2ydJqX/TlnEbEXIRlBYuBLgYoUGc37KNGEXirJRFe99jr4J0Bc3DpmxkfB+o
RDL+Q0q6ne+/rjgZcQW9nYF2wUu0Bh6VePFEM3l7fKcVbUfomAfMccEiS61obxTfCS8N+wSABJ3d
bbtJFOasgjOYNnKM14Gog13yMDcx35ln1CbC10fpSJywMXdHSnL83VmjQc+GcQJIz48wJu/Jh7DX
jPJaFvWtPiSy+i6TZFd0YgSRAdd2Q+uSHyOmtMhMoN+1NALI8aaKAE63Gz6v86ysev/c5E3z6K1w
gjO2JpO/SlWEv+NpzWodAk4cXiL80DbSWki4A6RfbRM4FMi7YsrhO5D2IXY9T4Yw3r493QSoSWFw
A57V3KyMuKZoGg/uxAOe4TzIXlii/2tmKLYh7Vlaf6lOX5EE4tw+e0wL/C6uaG+og/sG4xsP6tnw
/1HRmVO2C4EusmotD3LPu7w4gbVHs+U/Odg9FPO23jYlq5WsW0/W3OekQZS7R63feafySeXkRwNK
zIwCH16sUZRVbSRZG+QLtCD0m7IfCIXLbPSnZtb7H/cmCf5QkahnuCOp3CGz7tO6o3WlT2UY6Qjp
//xsO/qzl02ec3GHyr7I2e6Oh9GZp15LI9FDmWuJH6r51CA6sPQJWCSxRCdvZ72FqvqzQoeKfjQz
n46WSqfwzfYbrpatntuCKW2Zcx3Ymzly2YhN9yWoQgziCrPP8lqJVUt3P2Jz7HZO+yZAvQblCCGe
bvSUT966RAJZDLHwP4x1xlUiKXA0VnrtSBd3JmWA0ctneYWZlgjjObkuDc3a33+G7K0h7XPZBwmk
rZcTQuRsxrZxKYkx5tmHvWr9/lntv4mgkKK9IflNhQgfku4Pr/rfMFDH0GhNUHTl5Ss3j31xuj5q
rRKbZO86qg9+KmGevNhWzpkCUD+CGiFxEwTP7VfFFbmzLzORe3J1jqM5gn+dVJZ0uibSLXeoV7Et
kP0EPK1aRsyLVLfMF6z9VM/uErDfGVQmjeYAPOc5eGAAYuiBCOMjt+rkGKztC2QXg7/h9KEOLBNN
37MavjgRthx1sKsaLJWTQXJuOx8L1EQVRwLfnOy8ec3VulGTflDHAoQ1/5eFlviN7advSTWvhJz8
sH0GvT35wAvmHImkdqOzap71SYi9PflzRyqGzZM9POneGN//i2YoxigcShm17GOVbWLEAAu4REaD
WFulFYhO7XQT0HbGtnrr63HMfuuDKNT/iy+ARlgOzTL1nJ82cuX5KC2AUdvXokUh/t0xSaaubJOd
WihK9+rNzToheWzSExKXht4V/Wnla50qc+LarYtnFc7S00q5xyflJWZg7lh6a23Yd4BxEq8D7q1P
CgRgRGPPHTd4KCY9mgkwVQ4TCCzpxNZRSaNA7srpr7UZNxqjsFbEDhxG96Yy/0ClWpMCV5iB0Rrm
tjWwxFOjMssIU4Cj1/twdjaxY6jsFwFfY/acvBCxysj5iYMlwwl6F6+GVX5L+96lpabePu0jhdME
bNvSBlvlNB+PRreeelxwVyDZh9VRCaawFuXwtxk7/hcOVoaiO5WcQwHMHjW54uaNP0R3nW8hroEQ
oXrky1iurfp7ObH0gwVBC/QSVGhpXynRKF5W3jxQV4+BqFHsuLk1817pEYPHegXxcEU/+jHxzTR/
96UUtVEtkPlCb9nt4yH1YPBFsd/OAfgMxoV2cTP1l/D4l2LmAFm68QtMZJ9f949N6tDvjE5Crx69
ZcDc6CZQwnDaTOZxrp/zypdbIhRqjM+MjZJ8a46gIBBikdCaNdzV5weAYF8gYVhxzVAmK/O4Jhwa
9cc3erKJ1A5iMqt86nw2O1vYsNOuj1YxdBqVHN1oDvmPjbTVCYJIhj+gxbLDhurKv15YAHQfBIV/
CWEblBbVq+YK0BnTNOnlhlaxL4twmq7yxexkEJdXXAGv9uEwoA7Nrm6zJR2UDhxBdDJ3nfDLDBjt
/jHniWEpgCvadSLzK5Y7k/8CbatqwVn0LxH09Fm8fvrODMddUvbvoU7qHMT8eoSTS+IL/pLIInFr
Y2fQplytlK3qYl0SrKHYTObbvONlo/3H2sGBzeGkHYdc/6LaGoL+Oj4pV71x4lYeqj60QW9koISn
NtJTMNmGwQRtEv4s434Gav1jCufHKoCrKY3ucaAywa0+RWntjRABhsmLZDIjp8u6ZFdyr+COW3SX
6SP36W9quOgDtUdLmkBvvXlTjngWKjPIeyU10R9gtO1vRfzyXHWbEm9e6OcAxVzsWWW7kGHaVm9W
AVLhl7MD0q5HU7NH4CrD7sYldxMmHJJW/s4CJnH6/pKjX2DokQL83QUrIVUnRc3i1luk5WRmrYOv
WURDnJ5cIDSTLkWviX7EtYREIXFIdW+jeH7xSx3AKO7j88WAgwzCw8wBTtadjEhPme+gV7Stht0L
L90i5ciDJgujRjPP2HjUQIfBaAmMJt/0NGugPANBMDslF8a1o0XsTv4XmkRkx9N/uicPlIgGbI4E
gLq/ld9lEID9kuk4426jCxiUVkj71G2vBTu0Alm2s7Di4NIGD2CkgrOrYXXmuzi+0exci7f3Io6r
QBzARUIdRQoX3QLXIqpW0UbmvCIYaTtfrT0yvvyEW3QU5rPg3WvtzoisfvVSlODm3ASDzATHx3bj
a7ehAJRQAJ/8tDBucxUmo32Zyy+91+sOfyfvdQUjRaUCpIuK2Y8r5PdrstvMVnZ4nkaKp6BW0Wzu
nDYyNrE5Daxj9iSA5YasYKQbMYJIVYERJKTDoEzxgoaSz0wp0tdz2kTv80X2JJOyj5WGQh79+iXD
FewcYvLUEaFkqKfuqThUB9zUNTetbkNkrht0mdSUQj9SBoHOR3zd2qM9X9FBuWfIlGIz4Ww6TMF8
jZJq+q4ZQDZUG3x2kUcDquQ1VU1yB2X6cCavDCxuur2XlEx4Axp+jPyV4crscyDgQEu5AR5uhnIe
uYAD/83oU4FobRqOdVxIfU8jO94Cidi6jW/HLEja84gJuIskykXiNtg0h5DsKfIE3/ufyRdRqQ1u
z3Uak4569P0roRRlzw6UTPr2
`pragma protect end_protected

